`timescale 1ns / 1ps

module dct_8x8_stage_9_inner
(
    input wire clk,
    input wire rst,
    input wire [2048-1:0] i_data_in,
    input wire i_valid,
    output wire i_ready,
    output wire [2048-1:0] o_data_out,
    output wire o_valid,
    input wire o_ready
);

generate
/*
    Begin module dct_8x8_stage_9
*/
/*
    Wires declared by dct_8x8_stage_9
*/
wire FSM_dct_8x8_stage_9_0_in_ready;
wire FSM_dct_8x8_stage_9_0_out_valid;
/* End wires declared by dct_8x8_stage_9 */

/*
    Submodules of dct_8x8_stage_9
*/
reg [32-1:0] FSM_dct_8x8_stage_9_0_st_dummy_reg = 32'b0;

reg [32-1:0] FSM_dct_8x8_stage_9_0_t0;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t1;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t2;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t3;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t4;
reg [2048-1:0] FSM_dct_8x8_stage_9_0_t5;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t6;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t7;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t8;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t9;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t10;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t11;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t12;
reg [2048-1:0] FSM_dct_8x8_stage_9_0_t13;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t14;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t15;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t16;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t17;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t18;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t19;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t20;
reg [64-1:0] FSM_dct_8x8_stage_9_0_t21;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t22;
reg [2048-1:0] FSM_dct_8x8_stage_9_0_t23;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t24;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t25;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t26;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t27;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t28;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t29;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t30;
reg [2048-1:0] FSM_dct_8x8_stage_9_0_t31;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t32;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t33;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t34;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t35;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t36;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t37;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t38;
reg [64-1:0] FSM_dct_8x8_stage_9_0_t39;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t40;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t41;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t42;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t43;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t44;
reg [64-1:0] FSM_dct_8x8_stage_9_0_t45;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t46;
reg [2048-1:0] FSM_dct_8x8_stage_9_0_t47;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t48;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t49;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t50;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t51;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t52;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t53;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t54;
reg [64-1:0] FSM_dct_8x8_stage_9_0_t55;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t56;
reg [2048-1:0] FSM_dct_8x8_stage_9_0_t57;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t58;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t59;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t60;
reg [64-1:0] FSM_dct_8x8_stage_9_0_t61;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t62;
reg [2048-1:0] FSM_dct_8x8_stage_9_0_t63;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t64;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t65;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t66;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t67;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t68;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t69;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t70;
reg [2048-1:0] FSM_dct_8x8_stage_9_0_t71;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t72;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t73;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t74;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t75;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t76;
reg [2048-1:0] FSM_dct_8x8_stage_9_0_t77;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t78;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t79;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t80;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t81;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t82;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t83;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t84;
reg [2048-1:0] FSM_dct_8x8_stage_9_0_t85;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t86;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t87;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t88;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t89;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t90;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t91;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t92;
reg [64-1:0] FSM_dct_8x8_stage_9_0_t93;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t94;
reg [2048-1:0] FSM_dct_8x8_stage_9_0_t95;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t96;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t97;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t98;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t99;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t100;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t101;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t102;
reg [2048-1:0] FSM_dct_8x8_stage_9_0_t103;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t104;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t105;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t106;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t107;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t108;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t109;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t110;
reg [64-1:0] FSM_dct_8x8_stage_9_0_t111;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t112;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t113;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t114;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t115;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t116;
reg [64-1:0] FSM_dct_8x8_stage_9_0_t117;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t118;
reg [2048-1:0] FSM_dct_8x8_stage_9_0_t119;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t120;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t121;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t122;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t123;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t124;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t125;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t126;
reg [64-1:0] FSM_dct_8x8_stage_9_0_t127;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t128;
reg [2048-1:0] FSM_dct_8x8_stage_9_0_t129;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t130;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t131;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t132;
reg [64-1:0] FSM_dct_8x8_stage_9_0_t133;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t134;
reg [2048-1:0] FSM_dct_8x8_stage_9_0_t135;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t136;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t137;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t138;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t139;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t140;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t141;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t142;
reg [2048-1:0] FSM_dct_8x8_stage_9_0_t143;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t144;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t145;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t146;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t147;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t148;
reg [2048-1:0] FSM_dct_8x8_stage_9_0_t149;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t150;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t151;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t152;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t153;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t154;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t155;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t156;
reg [2048-1:0] FSM_dct_8x8_stage_9_0_t157;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t158;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t159;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t160;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t161;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t162;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t163;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t164;
reg [64-1:0] FSM_dct_8x8_stage_9_0_t165;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t166;
reg [2048-1:0] FSM_dct_8x8_stage_9_0_t167;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t168;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t169;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t170;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t171;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t172;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t173;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t174;
reg [2048-1:0] FSM_dct_8x8_stage_9_0_t175;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t176;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t177;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t178;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t179;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t180;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t181;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t182;
reg [64-1:0] FSM_dct_8x8_stage_9_0_t183;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t184;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t185;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t186;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t187;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t188;
reg [64-1:0] FSM_dct_8x8_stage_9_0_t189;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t190;
reg [2048-1:0] FSM_dct_8x8_stage_9_0_t191;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t192;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t193;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t194;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t195;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t196;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t197;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t198;
reg [64-1:0] FSM_dct_8x8_stage_9_0_t199;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t200;
reg [2048-1:0] FSM_dct_8x8_stage_9_0_t201;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t202;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t203;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t204;
reg [64-1:0] FSM_dct_8x8_stage_9_0_t205;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t206;
reg [2048-1:0] FSM_dct_8x8_stage_9_0_t207;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t208;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t209;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t210;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t211;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t212;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t213;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t214;
reg [2048-1:0] FSM_dct_8x8_stage_9_0_t215;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t216;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t217;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t218;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t219;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t220;
reg [2048-1:0] FSM_dct_8x8_stage_9_0_t221;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t222;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t223;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t224;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t225;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t226;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t227;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t228;
reg [2048-1:0] FSM_dct_8x8_stage_9_0_t229;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t230;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t231;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t232;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t233;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t234;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t235;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t236;
reg [64-1:0] FSM_dct_8x8_stage_9_0_t237;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t238;
reg [2048-1:0] FSM_dct_8x8_stage_9_0_t239;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t240;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t241;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t242;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t243;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t244;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t245;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t246;
reg [2048-1:0] FSM_dct_8x8_stage_9_0_t247;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t248;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t249;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t250;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t251;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t252;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t253;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t254;
reg [64-1:0] FSM_dct_8x8_stage_9_0_t255;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t256;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t257;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t258;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t259;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t260;
reg [64-1:0] FSM_dct_8x8_stage_9_0_t261;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t262;
reg [2048-1:0] FSM_dct_8x8_stage_9_0_t263;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t264;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t265;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t266;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t267;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t268;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t269;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t270;
reg [64-1:0] FSM_dct_8x8_stage_9_0_t271;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t272;
reg [2048-1:0] FSM_dct_8x8_stage_9_0_t273;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t274;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t275;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t276;
reg [64-1:0] FSM_dct_8x8_stage_9_0_t277;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t278;
reg [2048-1:0] FSM_dct_8x8_stage_9_0_t279;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t280;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t281;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t282;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t283;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t284;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t285;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t286;
reg [2048-1:0] FSM_dct_8x8_stage_9_0_t287;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t288;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t289;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t290;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t291;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t292;
reg [2048-1:0] FSM_dct_8x8_stage_9_0_t293;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t294;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t295;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t296;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t297;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t298;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t299;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t300;
reg [2048-1:0] FSM_dct_8x8_stage_9_0_t301;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t302;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t303;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t304;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t305;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t306;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t307;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t308;
reg [64-1:0] FSM_dct_8x8_stage_9_0_t309;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t310;
reg [2048-1:0] FSM_dct_8x8_stage_9_0_t311;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t312;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t313;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t314;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t315;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t316;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t317;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t318;
reg [2048-1:0] FSM_dct_8x8_stage_9_0_t319;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t320;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t321;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t322;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t323;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t324;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t325;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t326;
reg [64-1:0] FSM_dct_8x8_stage_9_0_t327;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t328;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t329;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t330;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t331;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t332;
reg [64-1:0] FSM_dct_8x8_stage_9_0_t333;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t334;
reg [2048-1:0] FSM_dct_8x8_stage_9_0_t335;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t336;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t337;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t338;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t339;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t340;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t341;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t342;
reg [64-1:0] FSM_dct_8x8_stage_9_0_t343;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t344;
reg [2048-1:0] FSM_dct_8x8_stage_9_0_t345;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t346;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t347;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t348;
reg [64-1:0] FSM_dct_8x8_stage_9_0_t349;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t350;
reg [2048-1:0] FSM_dct_8x8_stage_9_0_t351;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t352;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t353;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t354;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t355;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t356;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t357;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t358;
reg [2048-1:0] FSM_dct_8x8_stage_9_0_t359;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t360;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t361;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t362;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t363;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t364;
reg [2048-1:0] FSM_dct_8x8_stage_9_0_t365;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t366;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t367;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t368;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t369;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t370;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t371;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t372;
reg [2048-1:0] FSM_dct_8x8_stage_9_0_t373;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t374;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t375;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t376;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t377;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t378;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t379;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t380;
reg [64-1:0] FSM_dct_8x8_stage_9_0_t381;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t382;
reg [2048-1:0] FSM_dct_8x8_stage_9_0_t383;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t384;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t385;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t386;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t387;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t388;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t389;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t390;
reg [2048-1:0] FSM_dct_8x8_stage_9_0_t391;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t392;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t393;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t394;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t395;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t396;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t397;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t398;
reg [64-1:0] FSM_dct_8x8_stage_9_0_t399;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t400;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t401;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t402;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t403;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t404;
reg [64-1:0] FSM_dct_8x8_stage_9_0_t405;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t406;
reg [2048-1:0] FSM_dct_8x8_stage_9_0_t407;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t408;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t409;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t410;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t411;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t412;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t413;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t414;
reg [64-1:0] FSM_dct_8x8_stage_9_0_t415;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t416;
reg [2048-1:0] FSM_dct_8x8_stage_9_0_t417;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t418;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t419;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t420;
reg [64-1:0] FSM_dct_8x8_stage_9_0_t421;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t422;
reg [2048-1:0] FSM_dct_8x8_stage_9_0_t423;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t424;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t425;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t426;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t427;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t428;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t429;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t430;
reg [2048-1:0] FSM_dct_8x8_stage_9_0_t431;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t432;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t433;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t434;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t435;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t436;
reg [2048-1:0] FSM_dct_8x8_stage_9_0_t437;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t438;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t439;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t440;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t441;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t442;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t443;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t444;
reg [2048-1:0] FSM_dct_8x8_stage_9_0_t445;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t446;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t447;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t448;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t449;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t450;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t451;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t452;
reg [64-1:0] FSM_dct_8x8_stage_9_0_t453;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t454;
reg [2048-1:0] FSM_dct_8x8_stage_9_0_t455;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t456;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t457;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t458;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t459;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t460;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t461;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t462;
reg [2048-1:0] FSM_dct_8x8_stage_9_0_t463;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t464;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t465;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t466;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t467;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t468;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t469;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t470;
reg [64-1:0] FSM_dct_8x8_stage_9_0_t471;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t472;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t473;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t474;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t475;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t476;
reg [64-1:0] FSM_dct_8x8_stage_9_0_t477;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t478;
reg [2048-1:0] FSM_dct_8x8_stage_9_0_t479;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t480;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t481;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t482;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t483;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t484;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t485;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t486;
reg [64-1:0] FSM_dct_8x8_stage_9_0_t487;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t488;
reg [2048-1:0] FSM_dct_8x8_stage_9_0_t489;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t490;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t491;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t492;
reg [64-1:0] FSM_dct_8x8_stage_9_0_t493;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t494;
reg [2048-1:0] FSM_dct_8x8_stage_9_0_t495;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t496;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t497;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t498;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t499;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t500;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t501;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t502;
reg [2048-1:0] FSM_dct_8x8_stage_9_0_t503;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t504;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t505;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t506;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t507;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t508;
reg [2048-1:0] FSM_dct_8x8_stage_9_0_t509;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t510;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t511;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t512;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t513;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t514;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t515;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t516;
reg [2048-1:0] FSM_dct_8x8_stage_9_0_t517;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t518;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t519;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t520;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t521;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t522;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t523;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t524;
reg [64-1:0] FSM_dct_8x8_stage_9_0_t525;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t526;
reg [2048-1:0] FSM_dct_8x8_stage_9_0_t527;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t528;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t529;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t530;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t531;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t532;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t533;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t534;
reg [2048-1:0] FSM_dct_8x8_stage_9_0_t535;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t536;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t537;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t538;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t539;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t540;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t541;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t542;
reg [64-1:0] FSM_dct_8x8_stage_9_0_t543;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t544;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t545;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t546;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t547;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t548;
reg [64-1:0] FSM_dct_8x8_stage_9_0_t549;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t550;
reg [2048-1:0] FSM_dct_8x8_stage_9_0_t551;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t552;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t553;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t554;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t555;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t556;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t557;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t558;
reg [64-1:0] FSM_dct_8x8_stage_9_0_t559;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t560;
reg [2048-1:0] FSM_dct_8x8_stage_9_0_t561;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t562;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t563;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t564;
reg [64-1:0] FSM_dct_8x8_stage_9_0_t565;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t566;
reg [2048-1:0] FSM_dct_8x8_stage_9_0_t567;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t568;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t569;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t570;
reg [33-1:0] FSM_dct_8x8_stage_9_0_t571;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t572;
reg [6-1:0] FSM_dct_8x8_stage_9_0_t573;
reg [32-1:0] FSM_dct_8x8_stage_9_0_t574;
reg [2048-1:0] FSM_dct_8x8_stage_9_0_t575;

/*
    Wiring by dct_8x8_stage_9
*/
assign i_ready = FSM_dct_8x8_stage_9_0_in_ready;
assign o_data_out = FSM_dct_8x8_stage_9_0_t575;
assign o_valid = FSM_dct_8x8_stage_9_0_out_valid;
/* End wiring by dct_8x8_stage_9 */

assign FSM_dct_8x8_stage_9_0_out_valid = 1'b1;

initial begin
    FSM_dct_8x8_stage_9_0_t0 = 32'b0;
    FSM_dct_8x8_stage_9_0_t1 = FSM_dct_8x8_stage_9_0_t0[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t2 = 32'b0;
    FSM_dct_8x8_stage_9_0_t3 = FSM_dct_8x8_stage_9_0_t2[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t4 = i_data_in[FSM_dct_8x8_stage_9_0_t3 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t5 = 2048'b0;
    FSM_dct_8x8_stage_9_0_t5[FSM_dct_8x8_stage_9_0_t1 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t4;
    FSM_dct_8x8_stage_9_0_t6 = 32'b00000000000000000000000000001000 + 32'b0;
    FSM_dct_8x8_stage_9_0_t7 = FSM_dct_8x8_stage_9_0_t6[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t8 = FSM_dct_8x8_stage_9_0_t7[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t9 = 32'b00000000000000000000000000001000 + 32'b0;
    FSM_dct_8x8_stage_9_0_t10 = FSM_dct_8x8_stage_9_0_t9[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t11 = FSM_dct_8x8_stage_9_0_t10[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t12 = i_data_in[FSM_dct_8x8_stage_9_0_t11 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t13 = FSM_dct_8x8_stage_9_0_t5;
    FSM_dct_8x8_stage_9_0_t13[FSM_dct_8x8_stage_9_0_t8 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t12;
    FSM_dct_8x8_stage_9_0_t14 = 32'b00000000000000000000000000010000 + 32'b0;
    FSM_dct_8x8_stage_9_0_t15 = FSM_dct_8x8_stage_9_0_t14[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t16 = FSM_dct_8x8_stage_9_0_t15[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t17 = 32'b00000000000000000000000000010000 + 32'b0;
    FSM_dct_8x8_stage_9_0_t18 = FSM_dct_8x8_stage_9_0_t17[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t19 = FSM_dct_8x8_stage_9_0_t18[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t20 = i_data_in[FSM_dct_8x8_stage_9_0_t19 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t21 = FSM_dct_8x8_stage_9_0_t20 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t22 = FSM_dct_8x8_stage_9_0_t21[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t23 = FSM_dct_8x8_stage_9_0_t13;
    FSM_dct_8x8_stage_9_0_t23[FSM_dct_8x8_stage_9_0_t16 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t22;
    FSM_dct_8x8_stage_9_0_t24 = 32'b00000000000000000000000000011000 + 32'b0;
    FSM_dct_8x8_stage_9_0_t25 = FSM_dct_8x8_stage_9_0_t24[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t26 = FSM_dct_8x8_stage_9_0_t25[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t27 = 32'b00000000000000000000000000011000 + 32'b0;
    FSM_dct_8x8_stage_9_0_t28 = FSM_dct_8x8_stage_9_0_t27[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t29 = FSM_dct_8x8_stage_9_0_t28[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t30 = i_data_in[FSM_dct_8x8_stage_9_0_t29 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t31 = FSM_dct_8x8_stage_9_0_t23;
    FSM_dct_8x8_stage_9_0_t31[FSM_dct_8x8_stage_9_0_t26 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t30;
    FSM_dct_8x8_stage_9_0_t32 = 32'b00000000000000000000000000100000 + 32'b0;
    FSM_dct_8x8_stage_9_0_t33 = FSM_dct_8x8_stage_9_0_t32[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t34 = FSM_dct_8x8_stage_9_0_t33[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t35 = 32'b00000000000000000000000000100000 + 32'b0;
    FSM_dct_8x8_stage_9_0_t36 = FSM_dct_8x8_stage_9_0_t35[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t37 = FSM_dct_8x8_stage_9_0_t36[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t38 = i_data_in[FSM_dct_8x8_stage_9_0_t37 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t39 = FSM_dct_8x8_stage_9_0_t38 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t40 = FSM_dct_8x8_stage_9_0_t39[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t41 = 32'b00000000000000000000000000110000 + 32'b0;
    FSM_dct_8x8_stage_9_0_t42 = FSM_dct_8x8_stage_9_0_t41[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t43 = FSM_dct_8x8_stage_9_0_t42[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t44 = i_data_in[FSM_dct_8x8_stage_9_0_t43 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t45 = (FSM_dct_8x8_stage_9_0_t44 - FSM_dct_8x8_stage_9_0_t38) * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t46 = FSM_dct_8x8_stage_9_0_t45[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t47 = FSM_dct_8x8_stage_9_0_t31;
    FSM_dct_8x8_stage_9_0_t47[FSM_dct_8x8_stage_9_0_t34 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t40 - FSM_dct_8x8_stage_9_0_t46;
    FSM_dct_8x8_stage_9_0_t48 = 32'b00000000000000000000000000101000 + 32'b0;
    FSM_dct_8x8_stage_9_0_t49 = FSM_dct_8x8_stage_9_0_t48[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t50 = FSM_dct_8x8_stage_9_0_t49[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t51 = 32'b00000000000000000000000000101000 + 32'b0;
    FSM_dct_8x8_stage_9_0_t52 = FSM_dct_8x8_stage_9_0_t51[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t53 = FSM_dct_8x8_stage_9_0_t52[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t54 = i_data_in[FSM_dct_8x8_stage_9_0_t53 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t55 = FSM_dct_8x8_stage_9_0_t54 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t56 = FSM_dct_8x8_stage_9_0_t55[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t57 = FSM_dct_8x8_stage_9_0_t47;
    FSM_dct_8x8_stage_9_0_t57[FSM_dct_8x8_stage_9_0_t50 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t56;
    FSM_dct_8x8_stage_9_0_t58 = 32'b00000000000000000000000000110000 + 32'b0;
    FSM_dct_8x8_stage_9_0_t59 = FSM_dct_8x8_stage_9_0_t58[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t60 = FSM_dct_8x8_stage_9_0_t59[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t61 = FSM_dct_8x8_stage_9_0_t44 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t62 = FSM_dct_8x8_stage_9_0_t61[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t63 = FSM_dct_8x8_stage_9_0_t57;
    FSM_dct_8x8_stage_9_0_t63[FSM_dct_8x8_stage_9_0_t60 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t62 - FSM_dct_8x8_stage_9_0_t46;
    FSM_dct_8x8_stage_9_0_t64 = 32'b00000000000000000000000000111000 + 32'b0;
    FSM_dct_8x8_stage_9_0_t65 = FSM_dct_8x8_stage_9_0_t64[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t66 = FSM_dct_8x8_stage_9_0_t65[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t67 = 32'b00000000000000000000000000111000 + 32'b0;
    FSM_dct_8x8_stage_9_0_t68 = FSM_dct_8x8_stage_9_0_t67[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t69 = FSM_dct_8x8_stage_9_0_t68[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t70 = i_data_in[FSM_dct_8x8_stage_9_0_t69 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t71 = FSM_dct_8x8_stage_9_0_t63;
    FSM_dct_8x8_stage_9_0_t71[FSM_dct_8x8_stage_9_0_t66 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t70;
    FSM_dct_8x8_stage_9_0_t72 = 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_9_0_t73 = FSM_dct_8x8_stage_9_0_t72[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t74 = 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_9_0_t75 = FSM_dct_8x8_stage_9_0_t74[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t76 = i_data_in[FSM_dct_8x8_stage_9_0_t75 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t77 = FSM_dct_8x8_stage_9_0_t71;
    FSM_dct_8x8_stage_9_0_t77[FSM_dct_8x8_stage_9_0_t73 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t76;
    FSM_dct_8x8_stage_9_0_t78 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_9_0_t79 = FSM_dct_8x8_stage_9_0_t78[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t80 = FSM_dct_8x8_stage_9_0_t79[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t81 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_9_0_t82 = FSM_dct_8x8_stage_9_0_t81[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t83 = FSM_dct_8x8_stage_9_0_t82[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t84 = i_data_in[FSM_dct_8x8_stage_9_0_t83 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t85 = FSM_dct_8x8_stage_9_0_t77;
    FSM_dct_8x8_stage_9_0_t85[FSM_dct_8x8_stage_9_0_t80 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t84;
    FSM_dct_8x8_stage_9_0_t86 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_9_0_t87 = FSM_dct_8x8_stage_9_0_t86[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t88 = FSM_dct_8x8_stage_9_0_t87[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t89 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_9_0_t90 = FSM_dct_8x8_stage_9_0_t89[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t91 = FSM_dct_8x8_stage_9_0_t90[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t92 = i_data_in[FSM_dct_8x8_stage_9_0_t91 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t93 = FSM_dct_8x8_stage_9_0_t92 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t94 = FSM_dct_8x8_stage_9_0_t93[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t95 = FSM_dct_8x8_stage_9_0_t85;
    FSM_dct_8x8_stage_9_0_t95[FSM_dct_8x8_stage_9_0_t88 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t94;
    FSM_dct_8x8_stage_9_0_t96 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_9_0_t97 = FSM_dct_8x8_stage_9_0_t96[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t98 = FSM_dct_8x8_stage_9_0_t97[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t99 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_9_0_t100 = FSM_dct_8x8_stage_9_0_t99[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t101 = FSM_dct_8x8_stage_9_0_t100[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t102 = i_data_in[FSM_dct_8x8_stage_9_0_t101 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t103 = FSM_dct_8x8_stage_9_0_t95;
    FSM_dct_8x8_stage_9_0_t103[FSM_dct_8x8_stage_9_0_t98 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t102;
    FSM_dct_8x8_stage_9_0_t104 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_9_0_t105 = FSM_dct_8x8_stage_9_0_t104[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t106 = FSM_dct_8x8_stage_9_0_t105[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t107 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_9_0_t108 = FSM_dct_8x8_stage_9_0_t107[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t109 = FSM_dct_8x8_stage_9_0_t108[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t110 = i_data_in[FSM_dct_8x8_stage_9_0_t109 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t111 = FSM_dct_8x8_stage_9_0_t110 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t112 = FSM_dct_8x8_stage_9_0_t111[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t113 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_9_0_t114 = FSM_dct_8x8_stage_9_0_t113[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t115 = FSM_dct_8x8_stage_9_0_t114[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t116 = i_data_in[FSM_dct_8x8_stage_9_0_t115 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t117 = (FSM_dct_8x8_stage_9_0_t116 - FSM_dct_8x8_stage_9_0_t110) * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t118 = FSM_dct_8x8_stage_9_0_t117[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t119 = FSM_dct_8x8_stage_9_0_t103;
    FSM_dct_8x8_stage_9_0_t119[FSM_dct_8x8_stage_9_0_t106 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t112 - FSM_dct_8x8_stage_9_0_t118;
    FSM_dct_8x8_stage_9_0_t120 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_9_0_t121 = FSM_dct_8x8_stage_9_0_t120[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t122 = FSM_dct_8x8_stage_9_0_t121[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t123 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_9_0_t124 = FSM_dct_8x8_stage_9_0_t123[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t125 = FSM_dct_8x8_stage_9_0_t124[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t126 = i_data_in[FSM_dct_8x8_stage_9_0_t125 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t127 = FSM_dct_8x8_stage_9_0_t126 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t128 = FSM_dct_8x8_stage_9_0_t127[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t129 = FSM_dct_8x8_stage_9_0_t119;
    FSM_dct_8x8_stage_9_0_t129[FSM_dct_8x8_stage_9_0_t122 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t128;
    FSM_dct_8x8_stage_9_0_t130 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_9_0_t131 = FSM_dct_8x8_stage_9_0_t130[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t132 = FSM_dct_8x8_stage_9_0_t131[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t133 = FSM_dct_8x8_stage_9_0_t116 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t134 = FSM_dct_8x8_stage_9_0_t133[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t135 = FSM_dct_8x8_stage_9_0_t129;
    FSM_dct_8x8_stage_9_0_t135[FSM_dct_8x8_stage_9_0_t132 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t134 - FSM_dct_8x8_stage_9_0_t118;
    FSM_dct_8x8_stage_9_0_t136 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_9_0_t137 = FSM_dct_8x8_stage_9_0_t136[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t138 = FSM_dct_8x8_stage_9_0_t137[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t139 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_9_0_t140 = FSM_dct_8x8_stage_9_0_t139[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t141 = FSM_dct_8x8_stage_9_0_t140[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t142 = i_data_in[FSM_dct_8x8_stage_9_0_t141 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t143 = FSM_dct_8x8_stage_9_0_t135;
    FSM_dct_8x8_stage_9_0_t143[FSM_dct_8x8_stage_9_0_t138 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t142;
    FSM_dct_8x8_stage_9_0_t144 = 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_9_0_t145 = FSM_dct_8x8_stage_9_0_t144[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t146 = 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_9_0_t147 = FSM_dct_8x8_stage_9_0_t146[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t148 = i_data_in[FSM_dct_8x8_stage_9_0_t147 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t149 = FSM_dct_8x8_stage_9_0_t143;
    FSM_dct_8x8_stage_9_0_t149[FSM_dct_8x8_stage_9_0_t145 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t148;
    FSM_dct_8x8_stage_9_0_t150 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_9_0_t151 = FSM_dct_8x8_stage_9_0_t150[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t152 = FSM_dct_8x8_stage_9_0_t151[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t153 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_9_0_t154 = FSM_dct_8x8_stage_9_0_t153[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t155 = FSM_dct_8x8_stage_9_0_t154[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t156 = i_data_in[FSM_dct_8x8_stage_9_0_t155 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t157 = FSM_dct_8x8_stage_9_0_t149;
    FSM_dct_8x8_stage_9_0_t157[FSM_dct_8x8_stage_9_0_t152 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t156;
    FSM_dct_8x8_stage_9_0_t158 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_9_0_t159 = FSM_dct_8x8_stage_9_0_t158[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t160 = FSM_dct_8x8_stage_9_0_t159[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t161 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_9_0_t162 = FSM_dct_8x8_stage_9_0_t161[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t163 = FSM_dct_8x8_stage_9_0_t162[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t164 = i_data_in[FSM_dct_8x8_stage_9_0_t163 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t165 = FSM_dct_8x8_stage_9_0_t164 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t166 = FSM_dct_8x8_stage_9_0_t165[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t167 = FSM_dct_8x8_stage_9_0_t157;
    FSM_dct_8x8_stage_9_0_t167[FSM_dct_8x8_stage_9_0_t160 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t166;
    FSM_dct_8x8_stage_9_0_t168 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_9_0_t169 = FSM_dct_8x8_stage_9_0_t168[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t170 = FSM_dct_8x8_stage_9_0_t169[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t171 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_9_0_t172 = FSM_dct_8x8_stage_9_0_t171[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t173 = FSM_dct_8x8_stage_9_0_t172[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t174 = i_data_in[FSM_dct_8x8_stage_9_0_t173 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t175 = FSM_dct_8x8_stage_9_0_t167;
    FSM_dct_8x8_stage_9_0_t175[FSM_dct_8x8_stage_9_0_t170 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t174;
    FSM_dct_8x8_stage_9_0_t176 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_9_0_t177 = FSM_dct_8x8_stage_9_0_t176[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t178 = FSM_dct_8x8_stage_9_0_t177[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t179 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_9_0_t180 = FSM_dct_8x8_stage_9_0_t179[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t181 = FSM_dct_8x8_stage_9_0_t180[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t182 = i_data_in[FSM_dct_8x8_stage_9_0_t181 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t183 = FSM_dct_8x8_stage_9_0_t182 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t184 = FSM_dct_8x8_stage_9_0_t183[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t185 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_9_0_t186 = FSM_dct_8x8_stage_9_0_t185[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t187 = FSM_dct_8x8_stage_9_0_t186[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t188 = i_data_in[FSM_dct_8x8_stage_9_0_t187 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t189 = (FSM_dct_8x8_stage_9_0_t188 - FSM_dct_8x8_stage_9_0_t182) * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t190 = FSM_dct_8x8_stage_9_0_t189[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t191 = FSM_dct_8x8_stage_9_0_t175;
    FSM_dct_8x8_stage_9_0_t191[FSM_dct_8x8_stage_9_0_t178 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t184 - FSM_dct_8x8_stage_9_0_t190;
    FSM_dct_8x8_stage_9_0_t192 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_9_0_t193 = FSM_dct_8x8_stage_9_0_t192[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t194 = FSM_dct_8x8_stage_9_0_t193[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t195 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_9_0_t196 = FSM_dct_8x8_stage_9_0_t195[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t197 = FSM_dct_8x8_stage_9_0_t196[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t198 = i_data_in[FSM_dct_8x8_stage_9_0_t197 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t199 = FSM_dct_8x8_stage_9_0_t198 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t200 = FSM_dct_8x8_stage_9_0_t199[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t201 = FSM_dct_8x8_stage_9_0_t191;
    FSM_dct_8x8_stage_9_0_t201[FSM_dct_8x8_stage_9_0_t194 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t200;
    FSM_dct_8x8_stage_9_0_t202 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_9_0_t203 = FSM_dct_8x8_stage_9_0_t202[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t204 = FSM_dct_8x8_stage_9_0_t203[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t205 = FSM_dct_8x8_stage_9_0_t188 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t206 = FSM_dct_8x8_stage_9_0_t205[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t207 = FSM_dct_8x8_stage_9_0_t201;
    FSM_dct_8x8_stage_9_0_t207[FSM_dct_8x8_stage_9_0_t204 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t206 - FSM_dct_8x8_stage_9_0_t190;
    FSM_dct_8x8_stage_9_0_t208 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_9_0_t209 = FSM_dct_8x8_stage_9_0_t208[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t210 = FSM_dct_8x8_stage_9_0_t209[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t211 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_9_0_t212 = FSM_dct_8x8_stage_9_0_t211[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t213 = FSM_dct_8x8_stage_9_0_t212[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t214 = i_data_in[FSM_dct_8x8_stage_9_0_t213 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t215 = FSM_dct_8x8_stage_9_0_t207;
    FSM_dct_8x8_stage_9_0_t215[FSM_dct_8x8_stage_9_0_t210 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t214;
    FSM_dct_8x8_stage_9_0_t216 = 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_9_0_t217 = FSM_dct_8x8_stage_9_0_t216[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t218 = 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_9_0_t219 = FSM_dct_8x8_stage_9_0_t218[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t220 = i_data_in[FSM_dct_8x8_stage_9_0_t219 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t221 = FSM_dct_8x8_stage_9_0_t215;
    FSM_dct_8x8_stage_9_0_t221[FSM_dct_8x8_stage_9_0_t217 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t220;
    FSM_dct_8x8_stage_9_0_t222 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_9_0_t223 = FSM_dct_8x8_stage_9_0_t222[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t224 = FSM_dct_8x8_stage_9_0_t223[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t225 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_9_0_t226 = FSM_dct_8x8_stage_9_0_t225[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t227 = FSM_dct_8x8_stage_9_0_t226[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t228 = i_data_in[FSM_dct_8x8_stage_9_0_t227 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t229 = FSM_dct_8x8_stage_9_0_t221;
    FSM_dct_8x8_stage_9_0_t229[FSM_dct_8x8_stage_9_0_t224 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t228;
    FSM_dct_8x8_stage_9_0_t230 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_9_0_t231 = FSM_dct_8x8_stage_9_0_t230[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t232 = FSM_dct_8x8_stage_9_0_t231[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t233 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_9_0_t234 = FSM_dct_8x8_stage_9_0_t233[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t235 = FSM_dct_8x8_stage_9_0_t234[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t236 = i_data_in[FSM_dct_8x8_stage_9_0_t235 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t237 = FSM_dct_8x8_stage_9_0_t236 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t238 = FSM_dct_8x8_stage_9_0_t237[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t239 = FSM_dct_8x8_stage_9_0_t229;
    FSM_dct_8x8_stage_9_0_t239[FSM_dct_8x8_stage_9_0_t232 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t238;
    FSM_dct_8x8_stage_9_0_t240 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_9_0_t241 = FSM_dct_8x8_stage_9_0_t240[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t242 = FSM_dct_8x8_stage_9_0_t241[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t243 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_9_0_t244 = FSM_dct_8x8_stage_9_0_t243[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t245 = FSM_dct_8x8_stage_9_0_t244[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t246 = i_data_in[FSM_dct_8x8_stage_9_0_t245 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t247 = FSM_dct_8x8_stage_9_0_t239;
    FSM_dct_8x8_stage_9_0_t247[FSM_dct_8x8_stage_9_0_t242 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t246;
    FSM_dct_8x8_stage_9_0_t248 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_9_0_t249 = FSM_dct_8x8_stage_9_0_t248[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t250 = FSM_dct_8x8_stage_9_0_t249[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t251 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_9_0_t252 = FSM_dct_8x8_stage_9_0_t251[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t253 = FSM_dct_8x8_stage_9_0_t252[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t254 = i_data_in[FSM_dct_8x8_stage_9_0_t253 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t255 = FSM_dct_8x8_stage_9_0_t254 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t256 = FSM_dct_8x8_stage_9_0_t255[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t257 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_9_0_t258 = FSM_dct_8x8_stage_9_0_t257[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t259 = FSM_dct_8x8_stage_9_0_t258[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t260 = i_data_in[FSM_dct_8x8_stage_9_0_t259 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t261 = (FSM_dct_8x8_stage_9_0_t260 - FSM_dct_8x8_stage_9_0_t254) * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t262 = FSM_dct_8x8_stage_9_0_t261[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t263 = FSM_dct_8x8_stage_9_0_t247;
    FSM_dct_8x8_stage_9_0_t263[FSM_dct_8x8_stage_9_0_t250 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t256 - FSM_dct_8x8_stage_9_0_t262;
    FSM_dct_8x8_stage_9_0_t264 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_9_0_t265 = FSM_dct_8x8_stage_9_0_t264[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t266 = FSM_dct_8x8_stage_9_0_t265[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t267 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_9_0_t268 = FSM_dct_8x8_stage_9_0_t267[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t269 = FSM_dct_8x8_stage_9_0_t268[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t270 = i_data_in[FSM_dct_8x8_stage_9_0_t269 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t271 = FSM_dct_8x8_stage_9_0_t270 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t272 = FSM_dct_8x8_stage_9_0_t271[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t273 = FSM_dct_8x8_stage_9_0_t263;
    FSM_dct_8x8_stage_9_0_t273[FSM_dct_8x8_stage_9_0_t266 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t272;
    FSM_dct_8x8_stage_9_0_t274 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_9_0_t275 = FSM_dct_8x8_stage_9_0_t274[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t276 = FSM_dct_8x8_stage_9_0_t275[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t277 = FSM_dct_8x8_stage_9_0_t260 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t278 = FSM_dct_8x8_stage_9_0_t277[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t279 = FSM_dct_8x8_stage_9_0_t273;
    FSM_dct_8x8_stage_9_0_t279[FSM_dct_8x8_stage_9_0_t276 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t278 - FSM_dct_8x8_stage_9_0_t262;
    FSM_dct_8x8_stage_9_0_t280 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_9_0_t281 = FSM_dct_8x8_stage_9_0_t280[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t282 = FSM_dct_8x8_stage_9_0_t281[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t283 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_9_0_t284 = FSM_dct_8x8_stage_9_0_t283[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t285 = FSM_dct_8x8_stage_9_0_t284[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t286 = i_data_in[FSM_dct_8x8_stage_9_0_t285 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t287 = FSM_dct_8x8_stage_9_0_t279;
    FSM_dct_8x8_stage_9_0_t287[FSM_dct_8x8_stage_9_0_t282 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t286;
    FSM_dct_8x8_stage_9_0_t288 = 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_9_0_t289 = FSM_dct_8x8_stage_9_0_t288[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t290 = 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_9_0_t291 = FSM_dct_8x8_stage_9_0_t290[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t292 = i_data_in[FSM_dct_8x8_stage_9_0_t291 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t293 = FSM_dct_8x8_stage_9_0_t287;
    FSM_dct_8x8_stage_9_0_t293[FSM_dct_8x8_stage_9_0_t289 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t292;
    FSM_dct_8x8_stage_9_0_t294 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_9_0_t295 = FSM_dct_8x8_stage_9_0_t294[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t296 = FSM_dct_8x8_stage_9_0_t295[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t297 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_9_0_t298 = FSM_dct_8x8_stage_9_0_t297[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t299 = FSM_dct_8x8_stage_9_0_t298[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t300 = i_data_in[FSM_dct_8x8_stage_9_0_t299 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t301 = FSM_dct_8x8_stage_9_0_t293;
    FSM_dct_8x8_stage_9_0_t301[FSM_dct_8x8_stage_9_0_t296 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t300;
    FSM_dct_8x8_stage_9_0_t302 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_9_0_t303 = FSM_dct_8x8_stage_9_0_t302[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t304 = FSM_dct_8x8_stage_9_0_t303[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t305 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_9_0_t306 = FSM_dct_8x8_stage_9_0_t305[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t307 = FSM_dct_8x8_stage_9_0_t306[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t308 = i_data_in[FSM_dct_8x8_stage_9_0_t307 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t309 = FSM_dct_8x8_stage_9_0_t308 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t310 = FSM_dct_8x8_stage_9_0_t309[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t311 = FSM_dct_8x8_stage_9_0_t301;
    FSM_dct_8x8_stage_9_0_t311[FSM_dct_8x8_stage_9_0_t304 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t310;
    FSM_dct_8x8_stage_9_0_t312 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_9_0_t313 = FSM_dct_8x8_stage_9_0_t312[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t314 = FSM_dct_8x8_stage_9_0_t313[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t315 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_9_0_t316 = FSM_dct_8x8_stage_9_0_t315[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t317 = FSM_dct_8x8_stage_9_0_t316[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t318 = i_data_in[FSM_dct_8x8_stage_9_0_t317 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t319 = FSM_dct_8x8_stage_9_0_t311;
    FSM_dct_8x8_stage_9_0_t319[FSM_dct_8x8_stage_9_0_t314 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t318;
    FSM_dct_8x8_stage_9_0_t320 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_9_0_t321 = FSM_dct_8x8_stage_9_0_t320[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t322 = FSM_dct_8x8_stage_9_0_t321[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t323 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_9_0_t324 = FSM_dct_8x8_stage_9_0_t323[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t325 = FSM_dct_8x8_stage_9_0_t324[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t326 = i_data_in[FSM_dct_8x8_stage_9_0_t325 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t327 = FSM_dct_8x8_stage_9_0_t326 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t328 = FSM_dct_8x8_stage_9_0_t327[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t329 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_9_0_t330 = FSM_dct_8x8_stage_9_0_t329[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t331 = FSM_dct_8x8_stage_9_0_t330[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t332 = i_data_in[FSM_dct_8x8_stage_9_0_t331 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t333 = (FSM_dct_8x8_stage_9_0_t332 - FSM_dct_8x8_stage_9_0_t326) * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t334 = FSM_dct_8x8_stage_9_0_t333[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t335 = FSM_dct_8x8_stage_9_0_t319;
    FSM_dct_8x8_stage_9_0_t335[FSM_dct_8x8_stage_9_0_t322 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t328 - FSM_dct_8x8_stage_9_0_t334;
    FSM_dct_8x8_stage_9_0_t336 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_9_0_t337 = FSM_dct_8x8_stage_9_0_t336[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t338 = FSM_dct_8x8_stage_9_0_t337[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t339 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_9_0_t340 = FSM_dct_8x8_stage_9_0_t339[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t341 = FSM_dct_8x8_stage_9_0_t340[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t342 = i_data_in[FSM_dct_8x8_stage_9_0_t341 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t343 = FSM_dct_8x8_stage_9_0_t342 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t344 = FSM_dct_8x8_stage_9_0_t343[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t345 = FSM_dct_8x8_stage_9_0_t335;
    FSM_dct_8x8_stage_9_0_t345[FSM_dct_8x8_stage_9_0_t338 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t344;
    FSM_dct_8x8_stage_9_0_t346 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_9_0_t347 = FSM_dct_8x8_stage_9_0_t346[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t348 = FSM_dct_8x8_stage_9_0_t347[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t349 = FSM_dct_8x8_stage_9_0_t332 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t350 = FSM_dct_8x8_stage_9_0_t349[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t351 = FSM_dct_8x8_stage_9_0_t345;
    FSM_dct_8x8_stage_9_0_t351[FSM_dct_8x8_stage_9_0_t348 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t350 - FSM_dct_8x8_stage_9_0_t334;
    FSM_dct_8x8_stage_9_0_t352 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_9_0_t353 = FSM_dct_8x8_stage_9_0_t352[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t354 = FSM_dct_8x8_stage_9_0_t353[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t355 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_9_0_t356 = FSM_dct_8x8_stage_9_0_t355[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t357 = FSM_dct_8x8_stage_9_0_t356[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t358 = i_data_in[FSM_dct_8x8_stage_9_0_t357 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t359 = FSM_dct_8x8_stage_9_0_t351;
    FSM_dct_8x8_stage_9_0_t359[FSM_dct_8x8_stage_9_0_t354 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t358;
    FSM_dct_8x8_stage_9_0_t360 = 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_9_0_t361 = FSM_dct_8x8_stage_9_0_t360[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t362 = 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_9_0_t363 = FSM_dct_8x8_stage_9_0_t362[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t364 = i_data_in[FSM_dct_8x8_stage_9_0_t363 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t365 = FSM_dct_8x8_stage_9_0_t359;
    FSM_dct_8x8_stage_9_0_t365[FSM_dct_8x8_stage_9_0_t361 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t364;
    FSM_dct_8x8_stage_9_0_t366 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_9_0_t367 = FSM_dct_8x8_stage_9_0_t366[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t368 = FSM_dct_8x8_stage_9_0_t367[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t369 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_9_0_t370 = FSM_dct_8x8_stage_9_0_t369[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t371 = FSM_dct_8x8_stage_9_0_t370[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t372 = i_data_in[FSM_dct_8x8_stage_9_0_t371 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t373 = FSM_dct_8x8_stage_9_0_t365;
    FSM_dct_8x8_stage_9_0_t373[FSM_dct_8x8_stage_9_0_t368 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t372;
    FSM_dct_8x8_stage_9_0_t374 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_9_0_t375 = FSM_dct_8x8_stage_9_0_t374[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t376 = FSM_dct_8x8_stage_9_0_t375[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t377 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_9_0_t378 = FSM_dct_8x8_stage_9_0_t377[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t379 = FSM_dct_8x8_stage_9_0_t378[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t380 = i_data_in[FSM_dct_8x8_stage_9_0_t379 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t381 = FSM_dct_8x8_stage_9_0_t380 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t382 = FSM_dct_8x8_stage_9_0_t381[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t383 = FSM_dct_8x8_stage_9_0_t373;
    FSM_dct_8x8_stage_9_0_t383[FSM_dct_8x8_stage_9_0_t376 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t382;
    FSM_dct_8x8_stage_9_0_t384 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_9_0_t385 = FSM_dct_8x8_stage_9_0_t384[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t386 = FSM_dct_8x8_stage_9_0_t385[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t387 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_9_0_t388 = FSM_dct_8x8_stage_9_0_t387[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t389 = FSM_dct_8x8_stage_9_0_t388[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t390 = i_data_in[FSM_dct_8x8_stage_9_0_t389 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t391 = FSM_dct_8x8_stage_9_0_t383;
    FSM_dct_8x8_stage_9_0_t391[FSM_dct_8x8_stage_9_0_t386 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t390;
    FSM_dct_8x8_stage_9_0_t392 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_9_0_t393 = FSM_dct_8x8_stage_9_0_t392[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t394 = FSM_dct_8x8_stage_9_0_t393[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t395 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_9_0_t396 = FSM_dct_8x8_stage_9_0_t395[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t397 = FSM_dct_8x8_stage_9_0_t396[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t398 = i_data_in[FSM_dct_8x8_stage_9_0_t397 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t399 = FSM_dct_8x8_stage_9_0_t398 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t400 = FSM_dct_8x8_stage_9_0_t399[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t401 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_9_0_t402 = FSM_dct_8x8_stage_9_0_t401[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t403 = FSM_dct_8x8_stage_9_0_t402[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t404 = i_data_in[FSM_dct_8x8_stage_9_0_t403 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t405 = (FSM_dct_8x8_stage_9_0_t404 - FSM_dct_8x8_stage_9_0_t398) * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t406 = FSM_dct_8x8_stage_9_0_t405[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t407 = FSM_dct_8x8_stage_9_0_t391;
    FSM_dct_8x8_stage_9_0_t407[FSM_dct_8x8_stage_9_0_t394 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t400 - FSM_dct_8x8_stage_9_0_t406;
    FSM_dct_8x8_stage_9_0_t408 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_9_0_t409 = FSM_dct_8x8_stage_9_0_t408[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t410 = FSM_dct_8x8_stage_9_0_t409[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t411 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_9_0_t412 = FSM_dct_8x8_stage_9_0_t411[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t413 = FSM_dct_8x8_stage_9_0_t412[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t414 = i_data_in[FSM_dct_8x8_stage_9_0_t413 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t415 = FSM_dct_8x8_stage_9_0_t414 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t416 = FSM_dct_8x8_stage_9_0_t415[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t417 = FSM_dct_8x8_stage_9_0_t407;
    FSM_dct_8x8_stage_9_0_t417[FSM_dct_8x8_stage_9_0_t410 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t416;
    FSM_dct_8x8_stage_9_0_t418 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_9_0_t419 = FSM_dct_8x8_stage_9_0_t418[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t420 = FSM_dct_8x8_stage_9_0_t419[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t421 = FSM_dct_8x8_stage_9_0_t404 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t422 = FSM_dct_8x8_stage_9_0_t421[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t423 = FSM_dct_8x8_stage_9_0_t417;
    FSM_dct_8x8_stage_9_0_t423[FSM_dct_8x8_stage_9_0_t420 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t422 - FSM_dct_8x8_stage_9_0_t406;
    FSM_dct_8x8_stage_9_0_t424 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_9_0_t425 = FSM_dct_8x8_stage_9_0_t424[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t426 = FSM_dct_8x8_stage_9_0_t425[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t427 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_9_0_t428 = FSM_dct_8x8_stage_9_0_t427[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t429 = FSM_dct_8x8_stage_9_0_t428[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t430 = i_data_in[FSM_dct_8x8_stage_9_0_t429 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t431 = FSM_dct_8x8_stage_9_0_t423;
    FSM_dct_8x8_stage_9_0_t431[FSM_dct_8x8_stage_9_0_t426 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t430;
    FSM_dct_8x8_stage_9_0_t432 = 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_9_0_t433 = FSM_dct_8x8_stage_9_0_t432[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t434 = 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_9_0_t435 = FSM_dct_8x8_stage_9_0_t434[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t436 = i_data_in[FSM_dct_8x8_stage_9_0_t435 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t437 = FSM_dct_8x8_stage_9_0_t431;
    FSM_dct_8x8_stage_9_0_t437[FSM_dct_8x8_stage_9_0_t433 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t436;
    FSM_dct_8x8_stage_9_0_t438 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_9_0_t439 = FSM_dct_8x8_stage_9_0_t438[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t440 = FSM_dct_8x8_stage_9_0_t439[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t441 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_9_0_t442 = FSM_dct_8x8_stage_9_0_t441[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t443 = FSM_dct_8x8_stage_9_0_t442[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t444 = i_data_in[FSM_dct_8x8_stage_9_0_t443 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t445 = FSM_dct_8x8_stage_9_0_t437;
    FSM_dct_8x8_stage_9_0_t445[FSM_dct_8x8_stage_9_0_t440 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t444;
    FSM_dct_8x8_stage_9_0_t446 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_9_0_t447 = FSM_dct_8x8_stage_9_0_t446[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t448 = FSM_dct_8x8_stage_9_0_t447[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t449 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_9_0_t450 = FSM_dct_8x8_stage_9_0_t449[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t451 = FSM_dct_8x8_stage_9_0_t450[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t452 = i_data_in[FSM_dct_8x8_stage_9_0_t451 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t453 = FSM_dct_8x8_stage_9_0_t452 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t454 = FSM_dct_8x8_stage_9_0_t453[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t455 = FSM_dct_8x8_stage_9_0_t445;
    FSM_dct_8x8_stage_9_0_t455[FSM_dct_8x8_stage_9_0_t448 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t454;
    FSM_dct_8x8_stage_9_0_t456 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_9_0_t457 = FSM_dct_8x8_stage_9_0_t456[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t458 = FSM_dct_8x8_stage_9_0_t457[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t459 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_9_0_t460 = FSM_dct_8x8_stage_9_0_t459[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t461 = FSM_dct_8x8_stage_9_0_t460[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t462 = i_data_in[FSM_dct_8x8_stage_9_0_t461 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t463 = FSM_dct_8x8_stage_9_0_t455;
    FSM_dct_8x8_stage_9_0_t463[FSM_dct_8x8_stage_9_0_t458 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t462;
    FSM_dct_8x8_stage_9_0_t464 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_9_0_t465 = FSM_dct_8x8_stage_9_0_t464[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t466 = FSM_dct_8x8_stage_9_0_t465[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t467 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_9_0_t468 = FSM_dct_8x8_stage_9_0_t467[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t469 = FSM_dct_8x8_stage_9_0_t468[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t470 = i_data_in[FSM_dct_8x8_stage_9_0_t469 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t471 = FSM_dct_8x8_stage_9_0_t470 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t472 = FSM_dct_8x8_stage_9_0_t471[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t473 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_9_0_t474 = FSM_dct_8x8_stage_9_0_t473[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t475 = FSM_dct_8x8_stage_9_0_t474[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t476 = i_data_in[FSM_dct_8x8_stage_9_0_t475 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t477 = (FSM_dct_8x8_stage_9_0_t476 - FSM_dct_8x8_stage_9_0_t470) * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t478 = FSM_dct_8x8_stage_9_0_t477[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t479 = FSM_dct_8x8_stage_9_0_t463;
    FSM_dct_8x8_stage_9_0_t479[FSM_dct_8x8_stage_9_0_t466 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t472 - FSM_dct_8x8_stage_9_0_t478;
    FSM_dct_8x8_stage_9_0_t480 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_9_0_t481 = FSM_dct_8x8_stage_9_0_t480[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t482 = FSM_dct_8x8_stage_9_0_t481[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t483 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_9_0_t484 = FSM_dct_8x8_stage_9_0_t483[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t485 = FSM_dct_8x8_stage_9_0_t484[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t486 = i_data_in[FSM_dct_8x8_stage_9_0_t485 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t487 = FSM_dct_8x8_stage_9_0_t486 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t488 = FSM_dct_8x8_stage_9_0_t487[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t489 = FSM_dct_8x8_stage_9_0_t479;
    FSM_dct_8x8_stage_9_0_t489[FSM_dct_8x8_stage_9_0_t482 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t488;
    FSM_dct_8x8_stage_9_0_t490 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_9_0_t491 = FSM_dct_8x8_stage_9_0_t490[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t492 = FSM_dct_8x8_stage_9_0_t491[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t493 = FSM_dct_8x8_stage_9_0_t476 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t494 = FSM_dct_8x8_stage_9_0_t493[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t495 = FSM_dct_8x8_stage_9_0_t489;
    FSM_dct_8x8_stage_9_0_t495[FSM_dct_8x8_stage_9_0_t492 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t494 - FSM_dct_8x8_stage_9_0_t478;
    FSM_dct_8x8_stage_9_0_t496 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_9_0_t497 = FSM_dct_8x8_stage_9_0_t496[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t498 = FSM_dct_8x8_stage_9_0_t497[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t499 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_9_0_t500 = FSM_dct_8x8_stage_9_0_t499[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t501 = FSM_dct_8x8_stage_9_0_t500[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t502 = i_data_in[FSM_dct_8x8_stage_9_0_t501 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t503 = FSM_dct_8x8_stage_9_0_t495;
    FSM_dct_8x8_stage_9_0_t503[FSM_dct_8x8_stage_9_0_t498 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t502;
    FSM_dct_8x8_stage_9_0_t504 = 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_9_0_t505 = FSM_dct_8x8_stage_9_0_t504[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t506 = 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_9_0_t507 = FSM_dct_8x8_stage_9_0_t506[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t508 = i_data_in[FSM_dct_8x8_stage_9_0_t507 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t509 = FSM_dct_8x8_stage_9_0_t503;
    FSM_dct_8x8_stage_9_0_t509[FSM_dct_8x8_stage_9_0_t505 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t508;
    FSM_dct_8x8_stage_9_0_t510 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_9_0_t511 = FSM_dct_8x8_stage_9_0_t510[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t512 = FSM_dct_8x8_stage_9_0_t511[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t513 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_9_0_t514 = FSM_dct_8x8_stage_9_0_t513[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t515 = FSM_dct_8x8_stage_9_0_t514[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t516 = i_data_in[FSM_dct_8x8_stage_9_0_t515 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t517 = FSM_dct_8x8_stage_9_0_t509;
    FSM_dct_8x8_stage_9_0_t517[FSM_dct_8x8_stage_9_0_t512 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t516;
    FSM_dct_8x8_stage_9_0_t518 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_9_0_t519 = FSM_dct_8x8_stage_9_0_t518[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t520 = FSM_dct_8x8_stage_9_0_t519[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t521 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_9_0_t522 = FSM_dct_8x8_stage_9_0_t521[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t523 = FSM_dct_8x8_stage_9_0_t522[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t524 = i_data_in[FSM_dct_8x8_stage_9_0_t523 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t525 = FSM_dct_8x8_stage_9_0_t524 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t526 = FSM_dct_8x8_stage_9_0_t525[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t527 = FSM_dct_8x8_stage_9_0_t517;
    FSM_dct_8x8_stage_9_0_t527[FSM_dct_8x8_stage_9_0_t520 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t526;
    FSM_dct_8x8_stage_9_0_t528 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_9_0_t529 = FSM_dct_8x8_stage_9_0_t528[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t530 = FSM_dct_8x8_stage_9_0_t529[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t531 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_9_0_t532 = FSM_dct_8x8_stage_9_0_t531[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t533 = FSM_dct_8x8_stage_9_0_t532[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t534 = i_data_in[FSM_dct_8x8_stage_9_0_t533 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t535 = FSM_dct_8x8_stage_9_0_t527;
    FSM_dct_8x8_stage_9_0_t535[FSM_dct_8x8_stage_9_0_t530 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t534;
    FSM_dct_8x8_stage_9_0_t536 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_9_0_t537 = FSM_dct_8x8_stage_9_0_t536[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t538 = FSM_dct_8x8_stage_9_0_t537[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t539 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_9_0_t540 = FSM_dct_8x8_stage_9_0_t539[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t541 = FSM_dct_8x8_stage_9_0_t540[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t542 = i_data_in[FSM_dct_8x8_stage_9_0_t541 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t543 = FSM_dct_8x8_stage_9_0_t542 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t544 = FSM_dct_8x8_stage_9_0_t543[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t545 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_9_0_t546 = FSM_dct_8x8_stage_9_0_t545[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t547 = FSM_dct_8x8_stage_9_0_t546[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t548 = i_data_in[FSM_dct_8x8_stage_9_0_t547 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t549 = (FSM_dct_8x8_stage_9_0_t548 - FSM_dct_8x8_stage_9_0_t542) * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t550 = FSM_dct_8x8_stage_9_0_t549[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t551 = FSM_dct_8x8_stage_9_0_t535;
    FSM_dct_8x8_stage_9_0_t551[FSM_dct_8x8_stage_9_0_t538 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t544 - FSM_dct_8x8_stage_9_0_t550;
    FSM_dct_8x8_stage_9_0_t552 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_9_0_t553 = FSM_dct_8x8_stage_9_0_t552[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t554 = FSM_dct_8x8_stage_9_0_t553[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t555 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_9_0_t556 = FSM_dct_8x8_stage_9_0_t555[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t557 = FSM_dct_8x8_stage_9_0_t556[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t558 = i_data_in[FSM_dct_8x8_stage_9_0_t557 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t559 = FSM_dct_8x8_stage_9_0_t558 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t560 = FSM_dct_8x8_stage_9_0_t559[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t561 = FSM_dct_8x8_stage_9_0_t551;
    FSM_dct_8x8_stage_9_0_t561[FSM_dct_8x8_stage_9_0_t554 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t560;
    FSM_dct_8x8_stage_9_0_t562 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_9_0_t563 = FSM_dct_8x8_stage_9_0_t562[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t564 = FSM_dct_8x8_stage_9_0_t563[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t565 = FSM_dct_8x8_stage_9_0_t548 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t566 = FSM_dct_8x8_stage_9_0_t565[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t567 = FSM_dct_8x8_stage_9_0_t561;
    FSM_dct_8x8_stage_9_0_t567[FSM_dct_8x8_stage_9_0_t564 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t566 - FSM_dct_8x8_stage_9_0_t550;
    FSM_dct_8x8_stage_9_0_t568 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_9_0_t569 = FSM_dct_8x8_stage_9_0_t568[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t570 = FSM_dct_8x8_stage_9_0_t569[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t571 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_9_0_t572 = FSM_dct_8x8_stage_9_0_t571[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t573 = FSM_dct_8x8_stage_9_0_t572[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t574 = i_data_in[FSM_dct_8x8_stage_9_0_t573 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t575 = FSM_dct_8x8_stage_9_0_t567;
    FSM_dct_8x8_stage_9_0_t575[FSM_dct_8x8_stage_9_0_t570 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t574;
end

always @* begin
    FSM_dct_8x8_stage_9_0_t0 = 32'b0;
    FSM_dct_8x8_stage_9_0_t1 = FSM_dct_8x8_stage_9_0_t0[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t2 = 32'b0;
    FSM_dct_8x8_stage_9_0_t3 = FSM_dct_8x8_stage_9_0_t2[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t4 = i_data_in[FSM_dct_8x8_stage_9_0_t3 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t5 = 2048'b0;
    FSM_dct_8x8_stage_9_0_t5[FSM_dct_8x8_stage_9_0_t1 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t4;
    FSM_dct_8x8_stage_9_0_t6 = 32'b00000000000000000000000000001000 + 32'b0;
    FSM_dct_8x8_stage_9_0_t7 = FSM_dct_8x8_stage_9_0_t6[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t8 = FSM_dct_8x8_stage_9_0_t7[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t9 = 32'b00000000000000000000000000001000 + 32'b0;
    FSM_dct_8x8_stage_9_0_t10 = FSM_dct_8x8_stage_9_0_t9[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t11 = FSM_dct_8x8_stage_9_0_t10[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t12 = i_data_in[FSM_dct_8x8_stage_9_0_t11 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t13 = FSM_dct_8x8_stage_9_0_t5;
    FSM_dct_8x8_stage_9_0_t13[FSM_dct_8x8_stage_9_0_t8 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t12;
    FSM_dct_8x8_stage_9_0_t14 = 32'b00000000000000000000000000010000 + 32'b0;
    FSM_dct_8x8_stage_9_0_t15 = FSM_dct_8x8_stage_9_0_t14[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t16 = FSM_dct_8x8_stage_9_0_t15[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t17 = 32'b00000000000000000000000000010000 + 32'b0;
    FSM_dct_8x8_stage_9_0_t18 = FSM_dct_8x8_stage_9_0_t17[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t19 = FSM_dct_8x8_stage_9_0_t18[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t20 = i_data_in[FSM_dct_8x8_stage_9_0_t19 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t21 = FSM_dct_8x8_stage_9_0_t20 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t22 = FSM_dct_8x8_stage_9_0_t21[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t23 = FSM_dct_8x8_stage_9_0_t13;
    FSM_dct_8x8_stage_9_0_t23[FSM_dct_8x8_stage_9_0_t16 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t22;
    FSM_dct_8x8_stage_9_0_t24 = 32'b00000000000000000000000000011000 + 32'b0;
    FSM_dct_8x8_stage_9_0_t25 = FSM_dct_8x8_stage_9_0_t24[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t26 = FSM_dct_8x8_stage_9_0_t25[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t27 = 32'b00000000000000000000000000011000 + 32'b0;
    FSM_dct_8x8_stage_9_0_t28 = FSM_dct_8x8_stage_9_0_t27[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t29 = FSM_dct_8x8_stage_9_0_t28[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t30 = i_data_in[FSM_dct_8x8_stage_9_0_t29 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t31 = FSM_dct_8x8_stage_9_0_t23;
    FSM_dct_8x8_stage_9_0_t31[FSM_dct_8x8_stage_9_0_t26 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t30;
    FSM_dct_8x8_stage_9_0_t32 = 32'b00000000000000000000000000100000 + 32'b0;
    FSM_dct_8x8_stage_9_0_t33 = FSM_dct_8x8_stage_9_0_t32[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t34 = FSM_dct_8x8_stage_9_0_t33[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t35 = 32'b00000000000000000000000000100000 + 32'b0;
    FSM_dct_8x8_stage_9_0_t36 = FSM_dct_8x8_stage_9_0_t35[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t37 = FSM_dct_8x8_stage_9_0_t36[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t38 = i_data_in[FSM_dct_8x8_stage_9_0_t37 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t39 = FSM_dct_8x8_stage_9_0_t38 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t40 = FSM_dct_8x8_stage_9_0_t39[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t41 = 32'b00000000000000000000000000110000 + 32'b0;
    FSM_dct_8x8_stage_9_0_t42 = FSM_dct_8x8_stage_9_0_t41[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t43 = FSM_dct_8x8_stage_9_0_t42[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t44 = i_data_in[FSM_dct_8x8_stage_9_0_t43 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t45 = (FSM_dct_8x8_stage_9_0_t44 - FSM_dct_8x8_stage_9_0_t38) * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t46 = FSM_dct_8x8_stage_9_0_t45[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t47 = FSM_dct_8x8_stage_9_0_t31;
    FSM_dct_8x8_stage_9_0_t47[FSM_dct_8x8_stage_9_0_t34 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t40 - FSM_dct_8x8_stage_9_0_t46;
    FSM_dct_8x8_stage_9_0_t48 = 32'b00000000000000000000000000101000 + 32'b0;
    FSM_dct_8x8_stage_9_0_t49 = FSM_dct_8x8_stage_9_0_t48[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t50 = FSM_dct_8x8_stage_9_0_t49[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t51 = 32'b00000000000000000000000000101000 + 32'b0;
    FSM_dct_8x8_stage_9_0_t52 = FSM_dct_8x8_stage_9_0_t51[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t53 = FSM_dct_8x8_stage_9_0_t52[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t54 = i_data_in[FSM_dct_8x8_stage_9_0_t53 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t55 = FSM_dct_8x8_stage_9_0_t54 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t56 = FSM_dct_8x8_stage_9_0_t55[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t57 = FSM_dct_8x8_stage_9_0_t47;
    FSM_dct_8x8_stage_9_0_t57[FSM_dct_8x8_stage_9_0_t50 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t56;
    FSM_dct_8x8_stage_9_0_t58 = 32'b00000000000000000000000000110000 + 32'b0;
    FSM_dct_8x8_stage_9_0_t59 = FSM_dct_8x8_stage_9_0_t58[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t60 = FSM_dct_8x8_stage_9_0_t59[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t61 = FSM_dct_8x8_stage_9_0_t44 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t62 = FSM_dct_8x8_stage_9_0_t61[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t63 = FSM_dct_8x8_stage_9_0_t57;
    FSM_dct_8x8_stage_9_0_t63[FSM_dct_8x8_stage_9_0_t60 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t62 - FSM_dct_8x8_stage_9_0_t46;
    FSM_dct_8x8_stage_9_0_t64 = 32'b00000000000000000000000000111000 + 32'b0;
    FSM_dct_8x8_stage_9_0_t65 = FSM_dct_8x8_stage_9_0_t64[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t66 = FSM_dct_8x8_stage_9_0_t65[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t67 = 32'b00000000000000000000000000111000 + 32'b0;
    FSM_dct_8x8_stage_9_0_t68 = FSM_dct_8x8_stage_9_0_t67[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t69 = FSM_dct_8x8_stage_9_0_t68[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t70 = i_data_in[FSM_dct_8x8_stage_9_0_t69 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t71 = FSM_dct_8x8_stage_9_0_t63;
    FSM_dct_8x8_stage_9_0_t71[FSM_dct_8x8_stage_9_0_t66 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t70;
    FSM_dct_8x8_stage_9_0_t72 = 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_9_0_t73 = FSM_dct_8x8_stage_9_0_t72[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t74 = 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_9_0_t75 = FSM_dct_8x8_stage_9_0_t74[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t76 = i_data_in[FSM_dct_8x8_stage_9_0_t75 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t77 = FSM_dct_8x8_stage_9_0_t71;
    FSM_dct_8x8_stage_9_0_t77[FSM_dct_8x8_stage_9_0_t73 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t76;
    FSM_dct_8x8_stage_9_0_t78 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_9_0_t79 = FSM_dct_8x8_stage_9_0_t78[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t80 = FSM_dct_8x8_stage_9_0_t79[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t81 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_9_0_t82 = FSM_dct_8x8_stage_9_0_t81[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t83 = FSM_dct_8x8_stage_9_0_t82[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t84 = i_data_in[FSM_dct_8x8_stage_9_0_t83 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t85 = FSM_dct_8x8_stage_9_0_t77;
    FSM_dct_8x8_stage_9_0_t85[FSM_dct_8x8_stage_9_0_t80 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t84;
    FSM_dct_8x8_stage_9_0_t86 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_9_0_t87 = FSM_dct_8x8_stage_9_0_t86[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t88 = FSM_dct_8x8_stage_9_0_t87[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t89 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_9_0_t90 = FSM_dct_8x8_stage_9_0_t89[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t91 = FSM_dct_8x8_stage_9_0_t90[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t92 = i_data_in[FSM_dct_8x8_stage_9_0_t91 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t93 = FSM_dct_8x8_stage_9_0_t92 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t94 = FSM_dct_8x8_stage_9_0_t93[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t95 = FSM_dct_8x8_stage_9_0_t85;
    FSM_dct_8x8_stage_9_0_t95[FSM_dct_8x8_stage_9_0_t88 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t94;
    FSM_dct_8x8_stage_9_0_t96 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_9_0_t97 = FSM_dct_8x8_stage_9_0_t96[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t98 = FSM_dct_8x8_stage_9_0_t97[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t99 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_9_0_t100 = FSM_dct_8x8_stage_9_0_t99[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t101 = FSM_dct_8x8_stage_9_0_t100[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t102 = i_data_in[FSM_dct_8x8_stage_9_0_t101 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t103 = FSM_dct_8x8_stage_9_0_t95;
    FSM_dct_8x8_stage_9_0_t103[FSM_dct_8x8_stage_9_0_t98 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t102;
    FSM_dct_8x8_stage_9_0_t104 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_9_0_t105 = FSM_dct_8x8_stage_9_0_t104[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t106 = FSM_dct_8x8_stage_9_0_t105[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t107 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_9_0_t108 = FSM_dct_8x8_stage_9_0_t107[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t109 = FSM_dct_8x8_stage_9_0_t108[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t110 = i_data_in[FSM_dct_8x8_stage_9_0_t109 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t111 = FSM_dct_8x8_stage_9_0_t110 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t112 = FSM_dct_8x8_stage_9_0_t111[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t113 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_9_0_t114 = FSM_dct_8x8_stage_9_0_t113[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t115 = FSM_dct_8x8_stage_9_0_t114[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t116 = i_data_in[FSM_dct_8x8_stage_9_0_t115 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t117 = (FSM_dct_8x8_stage_9_0_t116 - FSM_dct_8x8_stage_9_0_t110) * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t118 = FSM_dct_8x8_stage_9_0_t117[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t119 = FSM_dct_8x8_stage_9_0_t103;
    FSM_dct_8x8_stage_9_0_t119[FSM_dct_8x8_stage_9_0_t106 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t112 - FSM_dct_8x8_stage_9_0_t118;
    FSM_dct_8x8_stage_9_0_t120 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_9_0_t121 = FSM_dct_8x8_stage_9_0_t120[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t122 = FSM_dct_8x8_stage_9_0_t121[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t123 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_9_0_t124 = FSM_dct_8x8_stage_9_0_t123[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t125 = FSM_dct_8x8_stage_9_0_t124[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t126 = i_data_in[FSM_dct_8x8_stage_9_0_t125 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t127 = FSM_dct_8x8_stage_9_0_t126 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t128 = FSM_dct_8x8_stage_9_0_t127[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t129 = FSM_dct_8x8_stage_9_0_t119;
    FSM_dct_8x8_stage_9_0_t129[FSM_dct_8x8_stage_9_0_t122 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t128;
    FSM_dct_8x8_stage_9_0_t130 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_9_0_t131 = FSM_dct_8x8_stage_9_0_t130[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t132 = FSM_dct_8x8_stage_9_0_t131[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t133 = FSM_dct_8x8_stage_9_0_t116 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t134 = FSM_dct_8x8_stage_9_0_t133[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t135 = FSM_dct_8x8_stage_9_0_t129;
    FSM_dct_8x8_stage_9_0_t135[FSM_dct_8x8_stage_9_0_t132 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t134 - FSM_dct_8x8_stage_9_0_t118;
    FSM_dct_8x8_stage_9_0_t136 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_9_0_t137 = FSM_dct_8x8_stage_9_0_t136[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t138 = FSM_dct_8x8_stage_9_0_t137[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t139 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_9_0_t140 = FSM_dct_8x8_stage_9_0_t139[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t141 = FSM_dct_8x8_stage_9_0_t140[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t142 = i_data_in[FSM_dct_8x8_stage_9_0_t141 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t143 = FSM_dct_8x8_stage_9_0_t135;
    FSM_dct_8x8_stage_9_0_t143[FSM_dct_8x8_stage_9_0_t138 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t142;
    FSM_dct_8x8_stage_9_0_t144 = 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_9_0_t145 = FSM_dct_8x8_stage_9_0_t144[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t146 = 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_9_0_t147 = FSM_dct_8x8_stage_9_0_t146[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t148 = i_data_in[FSM_dct_8x8_stage_9_0_t147 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t149 = FSM_dct_8x8_stage_9_0_t143;
    FSM_dct_8x8_stage_9_0_t149[FSM_dct_8x8_stage_9_0_t145 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t148;
    FSM_dct_8x8_stage_9_0_t150 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_9_0_t151 = FSM_dct_8x8_stage_9_0_t150[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t152 = FSM_dct_8x8_stage_9_0_t151[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t153 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_9_0_t154 = FSM_dct_8x8_stage_9_0_t153[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t155 = FSM_dct_8x8_stage_9_0_t154[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t156 = i_data_in[FSM_dct_8x8_stage_9_0_t155 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t157 = FSM_dct_8x8_stage_9_0_t149;
    FSM_dct_8x8_stage_9_0_t157[FSM_dct_8x8_stage_9_0_t152 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t156;
    FSM_dct_8x8_stage_9_0_t158 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_9_0_t159 = FSM_dct_8x8_stage_9_0_t158[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t160 = FSM_dct_8x8_stage_9_0_t159[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t161 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_9_0_t162 = FSM_dct_8x8_stage_9_0_t161[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t163 = FSM_dct_8x8_stage_9_0_t162[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t164 = i_data_in[FSM_dct_8x8_stage_9_0_t163 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t165 = FSM_dct_8x8_stage_9_0_t164 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t166 = FSM_dct_8x8_stage_9_0_t165[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t167 = FSM_dct_8x8_stage_9_0_t157;
    FSM_dct_8x8_stage_9_0_t167[FSM_dct_8x8_stage_9_0_t160 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t166;
    FSM_dct_8x8_stage_9_0_t168 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_9_0_t169 = FSM_dct_8x8_stage_9_0_t168[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t170 = FSM_dct_8x8_stage_9_0_t169[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t171 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_9_0_t172 = FSM_dct_8x8_stage_9_0_t171[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t173 = FSM_dct_8x8_stage_9_0_t172[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t174 = i_data_in[FSM_dct_8x8_stage_9_0_t173 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t175 = FSM_dct_8x8_stage_9_0_t167;
    FSM_dct_8x8_stage_9_0_t175[FSM_dct_8x8_stage_9_0_t170 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t174;
    FSM_dct_8x8_stage_9_0_t176 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_9_0_t177 = FSM_dct_8x8_stage_9_0_t176[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t178 = FSM_dct_8x8_stage_9_0_t177[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t179 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_9_0_t180 = FSM_dct_8x8_stage_9_0_t179[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t181 = FSM_dct_8x8_stage_9_0_t180[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t182 = i_data_in[FSM_dct_8x8_stage_9_0_t181 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t183 = FSM_dct_8x8_stage_9_0_t182 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t184 = FSM_dct_8x8_stage_9_0_t183[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t185 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_9_0_t186 = FSM_dct_8x8_stage_9_0_t185[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t187 = FSM_dct_8x8_stage_9_0_t186[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t188 = i_data_in[FSM_dct_8x8_stage_9_0_t187 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t189 = (FSM_dct_8x8_stage_9_0_t188 - FSM_dct_8x8_stage_9_0_t182) * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t190 = FSM_dct_8x8_stage_9_0_t189[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t191 = FSM_dct_8x8_stage_9_0_t175;
    FSM_dct_8x8_stage_9_0_t191[FSM_dct_8x8_stage_9_0_t178 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t184 - FSM_dct_8x8_stage_9_0_t190;
    FSM_dct_8x8_stage_9_0_t192 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_9_0_t193 = FSM_dct_8x8_stage_9_0_t192[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t194 = FSM_dct_8x8_stage_9_0_t193[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t195 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_9_0_t196 = FSM_dct_8x8_stage_9_0_t195[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t197 = FSM_dct_8x8_stage_9_0_t196[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t198 = i_data_in[FSM_dct_8x8_stage_9_0_t197 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t199 = FSM_dct_8x8_stage_9_0_t198 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t200 = FSM_dct_8x8_stage_9_0_t199[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t201 = FSM_dct_8x8_stage_9_0_t191;
    FSM_dct_8x8_stage_9_0_t201[FSM_dct_8x8_stage_9_0_t194 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t200;
    FSM_dct_8x8_stage_9_0_t202 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_9_0_t203 = FSM_dct_8x8_stage_9_0_t202[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t204 = FSM_dct_8x8_stage_9_0_t203[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t205 = FSM_dct_8x8_stage_9_0_t188 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t206 = FSM_dct_8x8_stage_9_0_t205[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t207 = FSM_dct_8x8_stage_9_0_t201;
    FSM_dct_8x8_stage_9_0_t207[FSM_dct_8x8_stage_9_0_t204 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t206 - FSM_dct_8x8_stage_9_0_t190;
    FSM_dct_8x8_stage_9_0_t208 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_9_0_t209 = FSM_dct_8x8_stage_9_0_t208[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t210 = FSM_dct_8x8_stage_9_0_t209[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t211 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_9_0_t212 = FSM_dct_8x8_stage_9_0_t211[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t213 = FSM_dct_8x8_stage_9_0_t212[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t214 = i_data_in[FSM_dct_8x8_stage_9_0_t213 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t215 = FSM_dct_8x8_stage_9_0_t207;
    FSM_dct_8x8_stage_9_0_t215[FSM_dct_8x8_stage_9_0_t210 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t214;
    FSM_dct_8x8_stage_9_0_t216 = 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_9_0_t217 = FSM_dct_8x8_stage_9_0_t216[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t218 = 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_9_0_t219 = FSM_dct_8x8_stage_9_0_t218[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t220 = i_data_in[FSM_dct_8x8_stage_9_0_t219 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t221 = FSM_dct_8x8_stage_9_0_t215;
    FSM_dct_8x8_stage_9_0_t221[FSM_dct_8x8_stage_9_0_t217 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t220;
    FSM_dct_8x8_stage_9_0_t222 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_9_0_t223 = FSM_dct_8x8_stage_9_0_t222[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t224 = FSM_dct_8x8_stage_9_0_t223[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t225 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_9_0_t226 = FSM_dct_8x8_stage_9_0_t225[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t227 = FSM_dct_8x8_stage_9_0_t226[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t228 = i_data_in[FSM_dct_8x8_stage_9_0_t227 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t229 = FSM_dct_8x8_stage_9_0_t221;
    FSM_dct_8x8_stage_9_0_t229[FSM_dct_8x8_stage_9_0_t224 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t228;
    FSM_dct_8x8_stage_9_0_t230 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_9_0_t231 = FSM_dct_8x8_stage_9_0_t230[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t232 = FSM_dct_8x8_stage_9_0_t231[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t233 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_9_0_t234 = FSM_dct_8x8_stage_9_0_t233[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t235 = FSM_dct_8x8_stage_9_0_t234[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t236 = i_data_in[FSM_dct_8x8_stage_9_0_t235 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t237 = FSM_dct_8x8_stage_9_0_t236 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t238 = FSM_dct_8x8_stage_9_0_t237[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t239 = FSM_dct_8x8_stage_9_0_t229;
    FSM_dct_8x8_stage_9_0_t239[FSM_dct_8x8_stage_9_0_t232 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t238;
    FSM_dct_8x8_stage_9_0_t240 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_9_0_t241 = FSM_dct_8x8_stage_9_0_t240[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t242 = FSM_dct_8x8_stage_9_0_t241[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t243 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_9_0_t244 = FSM_dct_8x8_stage_9_0_t243[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t245 = FSM_dct_8x8_stage_9_0_t244[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t246 = i_data_in[FSM_dct_8x8_stage_9_0_t245 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t247 = FSM_dct_8x8_stage_9_0_t239;
    FSM_dct_8x8_stage_9_0_t247[FSM_dct_8x8_stage_9_0_t242 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t246;
    FSM_dct_8x8_stage_9_0_t248 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_9_0_t249 = FSM_dct_8x8_stage_9_0_t248[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t250 = FSM_dct_8x8_stage_9_0_t249[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t251 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_9_0_t252 = FSM_dct_8x8_stage_9_0_t251[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t253 = FSM_dct_8x8_stage_9_0_t252[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t254 = i_data_in[FSM_dct_8x8_stage_9_0_t253 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t255 = FSM_dct_8x8_stage_9_0_t254 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t256 = FSM_dct_8x8_stage_9_0_t255[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t257 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_9_0_t258 = FSM_dct_8x8_stage_9_0_t257[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t259 = FSM_dct_8x8_stage_9_0_t258[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t260 = i_data_in[FSM_dct_8x8_stage_9_0_t259 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t261 = (FSM_dct_8x8_stage_9_0_t260 - FSM_dct_8x8_stage_9_0_t254) * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t262 = FSM_dct_8x8_stage_9_0_t261[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t263 = FSM_dct_8x8_stage_9_0_t247;
    FSM_dct_8x8_stage_9_0_t263[FSM_dct_8x8_stage_9_0_t250 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t256 - FSM_dct_8x8_stage_9_0_t262;
    FSM_dct_8x8_stage_9_0_t264 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_9_0_t265 = FSM_dct_8x8_stage_9_0_t264[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t266 = FSM_dct_8x8_stage_9_0_t265[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t267 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_9_0_t268 = FSM_dct_8x8_stage_9_0_t267[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t269 = FSM_dct_8x8_stage_9_0_t268[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t270 = i_data_in[FSM_dct_8x8_stage_9_0_t269 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t271 = FSM_dct_8x8_stage_9_0_t270 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t272 = FSM_dct_8x8_stage_9_0_t271[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t273 = FSM_dct_8x8_stage_9_0_t263;
    FSM_dct_8x8_stage_9_0_t273[FSM_dct_8x8_stage_9_0_t266 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t272;
    FSM_dct_8x8_stage_9_0_t274 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_9_0_t275 = FSM_dct_8x8_stage_9_0_t274[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t276 = FSM_dct_8x8_stage_9_0_t275[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t277 = FSM_dct_8x8_stage_9_0_t260 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t278 = FSM_dct_8x8_stage_9_0_t277[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t279 = FSM_dct_8x8_stage_9_0_t273;
    FSM_dct_8x8_stage_9_0_t279[FSM_dct_8x8_stage_9_0_t276 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t278 - FSM_dct_8x8_stage_9_0_t262;
    FSM_dct_8x8_stage_9_0_t280 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_9_0_t281 = FSM_dct_8x8_stage_9_0_t280[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t282 = FSM_dct_8x8_stage_9_0_t281[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t283 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_9_0_t284 = FSM_dct_8x8_stage_9_0_t283[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t285 = FSM_dct_8x8_stage_9_0_t284[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t286 = i_data_in[FSM_dct_8x8_stage_9_0_t285 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t287 = FSM_dct_8x8_stage_9_0_t279;
    FSM_dct_8x8_stage_9_0_t287[FSM_dct_8x8_stage_9_0_t282 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t286;
    FSM_dct_8x8_stage_9_0_t288 = 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_9_0_t289 = FSM_dct_8x8_stage_9_0_t288[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t290 = 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_9_0_t291 = FSM_dct_8x8_stage_9_0_t290[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t292 = i_data_in[FSM_dct_8x8_stage_9_0_t291 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t293 = FSM_dct_8x8_stage_9_0_t287;
    FSM_dct_8x8_stage_9_0_t293[FSM_dct_8x8_stage_9_0_t289 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t292;
    FSM_dct_8x8_stage_9_0_t294 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_9_0_t295 = FSM_dct_8x8_stage_9_0_t294[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t296 = FSM_dct_8x8_stage_9_0_t295[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t297 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_9_0_t298 = FSM_dct_8x8_stage_9_0_t297[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t299 = FSM_dct_8x8_stage_9_0_t298[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t300 = i_data_in[FSM_dct_8x8_stage_9_0_t299 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t301 = FSM_dct_8x8_stage_9_0_t293;
    FSM_dct_8x8_stage_9_0_t301[FSM_dct_8x8_stage_9_0_t296 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t300;
    FSM_dct_8x8_stage_9_0_t302 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_9_0_t303 = FSM_dct_8x8_stage_9_0_t302[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t304 = FSM_dct_8x8_stage_9_0_t303[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t305 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_9_0_t306 = FSM_dct_8x8_stage_9_0_t305[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t307 = FSM_dct_8x8_stage_9_0_t306[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t308 = i_data_in[FSM_dct_8x8_stage_9_0_t307 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t309 = FSM_dct_8x8_stage_9_0_t308 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t310 = FSM_dct_8x8_stage_9_0_t309[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t311 = FSM_dct_8x8_stage_9_0_t301;
    FSM_dct_8x8_stage_9_0_t311[FSM_dct_8x8_stage_9_0_t304 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t310;
    FSM_dct_8x8_stage_9_0_t312 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_9_0_t313 = FSM_dct_8x8_stage_9_0_t312[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t314 = FSM_dct_8x8_stage_9_0_t313[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t315 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_9_0_t316 = FSM_dct_8x8_stage_9_0_t315[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t317 = FSM_dct_8x8_stage_9_0_t316[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t318 = i_data_in[FSM_dct_8x8_stage_9_0_t317 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t319 = FSM_dct_8x8_stage_9_0_t311;
    FSM_dct_8x8_stage_9_0_t319[FSM_dct_8x8_stage_9_0_t314 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t318;
    FSM_dct_8x8_stage_9_0_t320 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_9_0_t321 = FSM_dct_8x8_stage_9_0_t320[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t322 = FSM_dct_8x8_stage_9_0_t321[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t323 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_9_0_t324 = FSM_dct_8x8_stage_9_0_t323[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t325 = FSM_dct_8x8_stage_9_0_t324[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t326 = i_data_in[FSM_dct_8x8_stage_9_0_t325 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t327 = FSM_dct_8x8_stage_9_0_t326 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t328 = FSM_dct_8x8_stage_9_0_t327[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t329 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_9_0_t330 = FSM_dct_8x8_stage_9_0_t329[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t331 = FSM_dct_8x8_stage_9_0_t330[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t332 = i_data_in[FSM_dct_8x8_stage_9_0_t331 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t333 = (FSM_dct_8x8_stage_9_0_t332 - FSM_dct_8x8_stage_9_0_t326) * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t334 = FSM_dct_8x8_stage_9_0_t333[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t335 = FSM_dct_8x8_stage_9_0_t319;
    FSM_dct_8x8_stage_9_0_t335[FSM_dct_8x8_stage_9_0_t322 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t328 - FSM_dct_8x8_stage_9_0_t334;
    FSM_dct_8x8_stage_9_0_t336 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_9_0_t337 = FSM_dct_8x8_stage_9_0_t336[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t338 = FSM_dct_8x8_stage_9_0_t337[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t339 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_9_0_t340 = FSM_dct_8x8_stage_9_0_t339[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t341 = FSM_dct_8x8_stage_9_0_t340[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t342 = i_data_in[FSM_dct_8x8_stage_9_0_t341 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t343 = FSM_dct_8x8_stage_9_0_t342 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t344 = FSM_dct_8x8_stage_9_0_t343[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t345 = FSM_dct_8x8_stage_9_0_t335;
    FSM_dct_8x8_stage_9_0_t345[FSM_dct_8x8_stage_9_0_t338 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t344;
    FSM_dct_8x8_stage_9_0_t346 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_9_0_t347 = FSM_dct_8x8_stage_9_0_t346[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t348 = FSM_dct_8x8_stage_9_0_t347[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t349 = FSM_dct_8x8_stage_9_0_t332 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t350 = FSM_dct_8x8_stage_9_0_t349[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t351 = FSM_dct_8x8_stage_9_0_t345;
    FSM_dct_8x8_stage_9_0_t351[FSM_dct_8x8_stage_9_0_t348 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t350 - FSM_dct_8x8_stage_9_0_t334;
    FSM_dct_8x8_stage_9_0_t352 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_9_0_t353 = FSM_dct_8x8_stage_9_0_t352[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t354 = FSM_dct_8x8_stage_9_0_t353[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t355 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_9_0_t356 = FSM_dct_8x8_stage_9_0_t355[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t357 = FSM_dct_8x8_stage_9_0_t356[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t358 = i_data_in[FSM_dct_8x8_stage_9_0_t357 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t359 = FSM_dct_8x8_stage_9_0_t351;
    FSM_dct_8x8_stage_9_0_t359[FSM_dct_8x8_stage_9_0_t354 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t358;
    FSM_dct_8x8_stage_9_0_t360 = 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_9_0_t361 = FSM_dct_8x8_stage_9_0_t360[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t362 = 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_9_0_t363 = FSM_dct_8x8_stage_9_0_t362[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t364 = i_data_in[FSM_dct_8x8_stage_9_0_t363 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t365 = FSM_dct_8x8_stage_9_0_t359;
    FSM_dct_8x8_stage_9_0_t365[FSM_dct_8x8_stage_9_0_t361 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t364;
    FSM_dct_8x8_stage_9_0_t366 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_9_0_t367 = FSM_dct_8x8_stage_9_0_t366[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t368 = FSM_dct_8x8_stage_9_0_t367[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t369 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_9_0_t370 = FSM_dct_8x8_stage_9_0_t369[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t371 = FSM_dct_8x8_stage_9_0_t370[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t372 = i_data_in[FSM_dct_8x8_stage_9_0_t371 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t373 = FSM_dct_8x8_stage_9_0_t365;
    FSM_dct_8x8_stage_9_0_t373[FSM_dct_8x8_stage_9_0_t368 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t372;
    FSM_dct_8x8_stage_9_0_t374 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_9_0_t375 = FSM_dct_8x8_stage_9_0_t374[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t376 = FSM_dct_8x8_stage_9_0_t375[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t377 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_9_0_t378 = FSM_dct_8x8_stage_9_0_t377[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t379 = FSM_dct_8x8_stage_9_0_t378[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t380 = i_data_in[FSM_dct_8x8_stage_9_0_t379 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t381 = FSM_dct_8x8_stage_9_0_t380 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t382 = FSM_dct_8x8_stage_9_0_t381[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t383 = FSM_dct_8x8_stage_9_0_t373;
    FSM_dct_8x8_stage_9_0_t383[FSM_dct_8x8_stage_9_0_t376 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t382;
    FSM_dct_8x8_stage_9_0_t384 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_9_0_t385 = FSM_dct_8x8_stage_9_0_t384[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t386 = FSM_dct_8x8_stage_9_0_t385[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t387 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_9_0_t388 = FSM_dct_8x8_stage_9_0_t387[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t389 = FSM_dct_8x8_stage_9_0_t388[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t390 = i_data_in[FSM_dct_8x8_stage_9_0_t389 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t391 = FSM_dct_8x8_stage_9_0_t383;
    FSM_dct_8x8_stage_9_0_t391[FSM_dct_8x8_stage_9_0_t386 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t390;
    FSM_dct_8x8_stage_9_0_t392 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_9_0_t393 = FSM_dct_8x8_stage_9_0_t392[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t394 = FSM_dct_8x8_stage_9_0_t393[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t395 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_9_0_t396 = FSM_dct_8x8_stage_9_0_t395[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t397 = FSM_dct_8x8_stage_9_0_t396[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t398 = i_data_in[FSM_dct_8x8_stage_9_0_t397 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t399 = FSM_dct_8x8_stage_9_0_t398 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t400 = FSM_dct_8x8_stage_9_0_t399[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t401 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_9_0_t402 = FSM_dct_8x8_stage_9_0_t401[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t403 = FSM_dct_8x8_stage_9_0_t402[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t404 = i_data_in[FSM_dct_8x8_stage_9_0_t403 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t405 = (FSM_dct_8x8_stage_9_0_t404 - FSM_dct_8x8_stage_9_0_t398) * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t406 = FSM_dct_8x8_stage_9_0_t405[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t407 = FSM_dct_8x8_stage_9_0_t391;
    FSM_dct_8x8_stage_9_0_t407[FSM_dct_8x8_stage_9_0_t394 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t400 - FSM_dct_8x8_stage_9_0_t406;
    FSM_dct_8x8_stage_9_0_t408 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_9_0_t409 = FSM_dct_8x8_stage_9_0_t408[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t410 = FSM_dct_8x8_stage_9_0_t409[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t411 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_9_0_t412 = FSM_dct_8x8_stage_9_0_t411[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t413 = FSM_dct_8x8_stage_9_0_t412[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t414 = i_data_in[FSM_dct_8x8_stage_9_0_t413 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t415 = FSM_dct_8x8_stage_9_0_t414 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t416 = FSM_dct_8x8_stage_9_0_t415[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t417 = FSM_dct_8x8_stage_9_0_t407;
    FSM_dct_8x8_stage_9_0_t417[FSM_dct_8x8_stage_9_0_t410 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t416;
    FSM_dct_8x8_stage_9_0_t418 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_9_0_t419 = FSM_dct_8x8_stage_9_0_t418[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t420 = FSM_dct_8x8_stage_9_0_t419[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t421 = FSM_dct_8x8_stage_9_0_t404 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t422 = FSM_dct_8x8_stage_9_0_t421[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t423 = FSM_dct_8x8_stage_9_0_t417;
    FSM_dct_8x8_stage_9_0_t423[FSM_dct_8x8_stage_9_0_t420 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t422 - FSM_dct_8x8_stage_9_0_t406;
    FSM_dct_8x8_stage_9_0_t424 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_9_0_t425 = FSM_dct_8x8_stage_9_0_t424[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t426 = FSM_dct_8x8_stage_9_0_t425[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t427 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_9_0_t428 = FSM_dct_8x8_stage_9_0_t427[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t429 = FSM_dct_8x8_stage_9_0_t428[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t430 = i_data_in[FSM_dct_8x8_stage_9_0_t429 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t431 = FSM_dct_8x8_stage_9_0_t423;
    FSM_dct_8x8_stage_9_0_t431[FSM_dct_8x8_stage_9_0_t426 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t430;
    FSM_dct_8x8_stage_9_0_t432 = 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_9_0_t433 = FSM_dct_8x8_stage_9_0_t432[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t434 = 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_9_0_t435 = FSM_dct_8x8_stage_9_0_t434[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t436 = i_data_in[FSM_dct_8x8_stage_9_0_t435 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t437 = FSM_dct_8x8_stage_9_0_t431;
    FSM_dct_8x8_stage_9_0_t437[FSM_dct_8x8_stage_9_0_t433 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t436;
    FSM_dct_8x8_stage_9_0_t438 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_9_0_t439 = FSM_dct_8x8_stage_9_0_t438[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t440 = FSM_dct_8x8_stage_9_0_t439[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t441 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_9_0_t442 = FSM_dct_8x8_stage_9_0_t441[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t443 = FSM_dct_8x8_stage_9_0_t442[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t444 = i_data_in[FSM_dct_8x8_stage_9_0_t443 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t445 = FSM_dct_8x8_stage_9_0_t437;
    FSM_dct_8x8_stage_9_0_t445[FSM_dct_8x8_stage_9_0_t440 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t444;
    FSM_dct_8x8_stage_9_0_t446 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_9_0_t447 = FSM_dct_8x8_stage_9_0_t446[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t448 = FSM_dct_8x8_stage_9_0_t447[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t449 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_9_0_t450 = FSM_dct_8x8_stage_9_0_t449[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t451 = FSM_dct_8x8_stage_9_0_t450[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t452 = i_data_in[FSM_dct_8x8_stage_9_0_t451 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t453 = FSM_dct_8x8_stage_9_0_t452 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t454 = FSM_dct_8x8_stage_9_0_t453[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t455 = FSM_dct_8x8_stage_9_0_t445;
    FSM_dct_8x8_stage_9_0_t455[FSM_dct_8x8_stage_9_0_t448 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t454;
    FSM_dct_8x8_stage_9_0_t456 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_9_0_t457 = FSM_dct_8x8_stage_9_0_t456[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t458 = FSM_dct_8x8_stage_9_0_t457[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t459 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_9_0_t460 = FSM_dct_8x8_stage_9_0_t459[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t461 = FSM_dct_8x8_stage_9_0_t460[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t462 = i_data_in[FSM_dct_8x8_stage_9_0_t461 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t463 = FSM_dct_8x8_stage_9_0_t455;
    FSM_dct_8x8_stage_9_0_t463[FSM_dct_8x8_stage_9_0_t458 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t462;
    FSM_dct_8x8_stage_9_0_t464 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_9_0_t465 = FSM_dct_8x8_stage_9_0_t464[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t466 = FSM_dct_8x8_stage_9_0_t465[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t467 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_9_0_t468 = FSM_dct_8x8_stage_9_0_t467[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t469 = FSM_dct_8x8_stage_9_0_t468[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t470 = i_data_in[FSM_dct_8x8_stage_9_0_t469 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t471 = FSM_dct_8x8_stage_9_0_t470 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t472 = FSM_dct_8x8_stage_9_0_t471[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t473 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_9_0_t474 = FSM_dct_8x8_stage_9_0_t473[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t475 = FSM_dct_8x8_stage_9_0_t474[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t476 = i_data_in[FSM_dct_8x8_stage_9_0_t475 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t477 = (FSM_dct_8x8_stage_9_0_t476 - FSM_dct_8x8_stage_9_0_t470) * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t478 = FSM_dct_8x8_stage_9_0_t477[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t479 = FSM_dct_8x8_stage_9_0_t463;
    FSM_dct_8x8_stage_9_0_t479[FSM_dct_8x8_stage_9_0_t466 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t472 - FSM_dct_8x8_stage_9_0_t478;
    FSM_dct_8x8_stage_9_0_t480 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_9_0_t481 = FSM_dct_8x8_stage_9_0_t480[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t482 = FSM_dct_8x8_stage_9_0_t481[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t483 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_9_0_t484 = FSM_dct_8x8_stage_9_0_t483[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t485 = FSM_dct_8x8_stage_9_0_t484[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t486 = i_data_in[FSM_dct_8x8_stage_9_0_t485 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t487 = FSM_dct_8x8_stage_9_0_t486 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t488 = FSM_dct_8x8_stage_9_0_t487[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t489 = FSM_dct_8x8_stage_9_0_t479;
    FSM_dct_8x8_stage_9_0_t489[FSM_dct_8x8_stage_9_0_t482 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t488;
    FSM_dct_8x8_stage_9_0_t490 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_9_0_t491 = FSM_dct_8x8_stage_9_0_t490[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t492 = FSM_dct_8x8_stage_9_0_t491[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t493 = FSM_dct_8x8_stage_9_0_t476 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t494 = FSM_dct_8x8_stage_9_0_t493[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t495 = FSM_dct_8x8_stage_9_0_t489;
    FSM_dct_8x8_stage_9_0_t495[FSM_dct_8x8_stage_9_0_t492 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t494 - FSM_dct_8x8_stage_9_0_t478;
    FSM_dct_8x8_stage_9_0_t496 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_9_0_t497 = FSM_dct_8x8_stage_9_0_t496[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t498 = FSM_dct_8x8_stage_9_0_t497[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t499 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_9_0_t500 = FSM_dct_8x8_stage_9_0_t499[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t501 = FSM_dct_8x8_stage_9_0_t500[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t502 = i_data_in[FSM_dct_8x8_stage_9_0_t501 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t503 = FSM_dct_8x8_stage_9_0_t495;
    FSM_dct_8x8_stage_9_0_t503[FSM_dct_8x8_stage_9_0_t498 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t502;
    FSM_dct_8x8_stage_9_0_t504 = 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_9_0_t505 = FSM_dct_8x8_stage_9_0_t504[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t506 = 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_9_0_t507 = FSM_dct_8x8_stage_9_0_t506[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t508 = i_data_in[FSM_dct_8x8_stage_9_0_t507 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t509 = FSM_dct_8x8_stage_9_0_t503;
    FSM_dct_8x8_stage_9_0_t509[FSM_dct_8x8_stage_9_0_t505 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t508;
    FSM_dct_8x8_stage_9_0_t510 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_9_0_t511 = FSM_dct_8x8_stage_9_0_t510[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t512 = FSM_dct_8x8_stage_9_0_t511[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t513 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_9_0_t514 = FSM_dct_8x8_stage_9_0_t513[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t515 = FSM_dct_8x8_stage_9_0_t514[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t516 = i_data_in[FSM_dct_8x8_stage_9_0_t515 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t517 = FSM_dct_8x8_stage_9_0_t509;
    FSM_dct_8x8_stage_9_0_t517[FSM_dct_8x8_stage_9_0_t512 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t516;
    FSM_dct_8x8_stage_9_0_t518 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_9_0_t519 = FSM_dct_8x8_stage_9_0_t518[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t520 = FSM_dct_8x8_stage_9_0_t519[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t521 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_9_0_t522 = FSM_dct_8x8_stage_9_0_t521[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t523 = FSM_dct_8x8_stage_9_0_t522[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t524 = i_data_in[FSM_dct_8x8_stage_9_0_t523 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t525 = FSM_dct_8x8_stage_9_0_t524 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t526 = FSM_dct_8x8_stage_9_0_t525[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t527 = FSM_dct_8x8_stage_9_0_t517;
    FSM_dct_8x8_stage_9_0_t527[FSM_dct_8x8_stage_9_0_t520 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t526;
    FSM_dct_8x8_stage_9_0_t528 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_9_0_t529 = FSM_dct_8x8_stage_9_0_t528[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t530 = FSM_dct_8x8_stage_9_0_t529[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t531 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_9_0_t532 = FSM_dct_8x8_stage_9_0_t531[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t533 = FSM_dct_8x8_stage_9_0_t532[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t534 = i_data_in[FSM_dct_8x8_stage_9_0_t533 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t535 = FSM_dct_8x8_stage_9_0_t527;
    FSM_dct_8x8_stage_9_0_t535[FSM_dct_8x8_stage_9_0_t530 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t534;
    FSM_dct_8x8_stage_9_0_t536 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_9_0_t537 = FSM_dct_8x8_stage_9_0_t536[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t538 = FSM_dct_8x8_stage_9_0_t537[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t539 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_9_0_t540 = FSM_dct_8x8_stage_9_0_t539[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t541 = FSM_dct_8x8_stage_9_0_t540[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t542 = i_data_in[FSM_dct_8x8_stage_9_0_t541 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t543 = FSM_dct_8x8_stage_9_0_t542 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t544 = FSM_dct_8x8_stage_9_0_t543[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t545 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_9_0_t546 = FSM_dct_8x8_stage_9_0_t545[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t547 = FSM_dct_8x8_stage_9_0_t546[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t548 = i_data_in[FSM_dct_8x8_stage_9_0_t547 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t549 = (FSM_dct_8x8_stage_9_0_t548 - FSM_dct_8x8_stage_9_0_t542) * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t550 = FSM_dct_8x8_stage_9_0_t549[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t551 = FSM_dct_8x8_stage_9_0_t535;
    FSM_dct_8x8_stage_9_0_t551[FSM_dct_8x8_stage_9_0_t538 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t544 - FSM_dct_8x8_stage_9_0_t550;
    FSM_dct_8x8_stage_9_0_t552 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_9_0_t553 = FSM_dct_8x8_stage_9_0_t552[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t554 = FSM_dct_8x8_stage_9_0_t553[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t555 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_9_0_t556 = FSM_dct_8x8_stage_9_0_t555[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t557 = FSM_dct_8x8_stage_9_0_t556[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t558 = i_data_in[FSM_dct_8x8_stage_9_0_t557 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t559 = FSM_dct_8x8_stage_9_0_t558 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t560 = FSM_dct_8x8_stage_9_0_t559[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t561 = FSM_dct_8x8_stage_9_0_t551;
    FSM_dct_8x8_stage_9_0_t561[FSM_dct_8x8_stage_9_0_t554 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t560;
    FSM_dct_8x8_stage_9_0_t562 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_9_0_t563 = FSM_dct_8x8_stage_9_0_t562[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t564 = FSM_dct_8x8_stage_9_0_t563[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t565 = FSM_dct_8x8_stage_9_0_t548 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_9_0_t566 = FSM_dct_8x8_stage_9_0_t565[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t567 = FSM_dct_8x8_stage_9_0_t561;
    FSM_dct_8x8_stage_9_0_t567[FSM_dct_8x8_stage_9_0_t564 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t566 - FSM_dct_8x8_stage_9_0_t550;
    FSM_dct_8x8_stage_9_0_t568 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_9_0_t569 = FSM_dct_8x8_stage_9_0_t568[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t570 = FSM_dct_8x8_stage_9_0_t569[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t571 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_9_0_t572 = FSM_dct_8x8_stage_9_0_t571[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_9_0_t573 = FSM_dct_8x8_stage_9_0_t572[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_9_0_t574 = i_data_in[FSM_dct_8x8_stage_9_0_t573 * 32 +: 32];
    FSM_dct_8x8_stage_9_0_t575 = FSM_dct_8x8_stage_9_0_t567;
    FSM_dct_8x8_stage_9_0_t575[FSM_dct_8x8_stage_9_0_t570 * 32 +: 32] = FSM_dct_8x8_stage_9_0_t574;
end

assign FSM_dct_8x8_stage_9_0_in_ready = 1'b1;

always @(posedge clk) begin
    FSM_dct_8x8_stage_9_0_st_dummy_reg <= FSM_dct_8x8_stage_9_0_st_dummy_reg;
    if (rst) begin
        FSM_dct_8x8_stage_9_0_st_dummy_reg <= 32'b0;
    end
end
/* End submodules of dct_8x8_stage_9 */
/* End module dct_8x8_stage_9 */
endgenerate
endmodule
