`timescale 1ns / 1ps

module sub_bytes_inner
(
    input wire clk,
    input wire rst,
    input wire [64-1:0] i_higher_bits,
    input wire [64-1:0] i_lower_bits,
    input wire i_valid,
    output wire i_ready,
    output wire [64-1:0] o_higher_out,
    output wire [64-1:0] o_lower_out,
    output wire o_valid,
    input wire o_ready
);

generate
/*
    Begin module sub_bytes
*/
/*
    Wires declared by sub_bytes
*/
wire FSM_sub_bytes_0_in_ready;
wire [64-1:0] FSM_sub_bytes_0_out_higher_out;
wire [64-1:0] FSM_sub_bytes_0_out_lower_out;
wire FSM_sub_bytes_0_out_valid;
/* End wires declared by sub_bytes */

/*
    Submodules of sub_bytes
*/
reg [64-1:0] FSM_sub_bytes_0_st_dummy_reg = 64'b0;

reg [1024-1:0] FSM_sub_bytes_0_t0;
reg [64-1:0] FSM_sub_bytes_0_t1;
reg [6-1:0] FSM_sub_bytes_0_t2;
reg [64-1:0] FSM_sub_bytes_0_t3;
reg [6-1:0] FSM_sub_bytes_0_t4;
reg [64-1:0] FSM_sub_bytes_0_t5;
reg [6-1:0] FSM_sub_bytes_0_t6;
reg [64-1:0] FSM_sub_bytes_0_t7;
reg [6-1:0] FSM_sub_bytes_0_t8;
reg [64-1:0] FSM_sub_bytes_0_t9;
reg [6-1:0] FSM_sub_bytes_0_t10;
reg [64-1:0] FSM_sub_bytes_0_t11;
reg [6-1:0] FSM_sub_bytes_0_t12;
reg [64-1:0] FSM_sub_bytes_0_t13;
reg [6-1:0] FSM_sub_bytes_0_t14;
reg [64-1:0] FSM_sub_bytes_0_t15;
reg [6-1:0] FSM_sub_bytes_0_t16;
reg [64-1:0] FSM_sub_bytes_0_t17;
reg [6-1:0] FSM_sub_bytes_0_t18;
reg [64-1:0] FSM_sub_bytes_0_t19;
reg [6-1:0] FSM_sub_bytes_0_t20;
reg [64-1:0] FSM_sub_bytes_0_t21;
reg [6-1:0] FSM_sub_bytes_0_t22;
reg [64-1:0] FSM_sub_bytes_0_t23;
reg [6-1:0] FSM_sub_bytes_0_t24;
reg [64-1:0] FSM_sub_bytes_0_t25;
reg [6-1:0] FSM_sub_bytes_0_t26;
reg [64-1:0] FSM_sub_bytes_0_t27;
reg [6-1:0] FSM_sub_bytes_0_t28;
reg [64-1:0] FSM_sub_bytes_0_t29;
reg [4-1:0] FSM_sub_bytes_0_t30;
reg [16384-1:0] FSM_sub_bytes_0_t31;
reg [64-1:0] FSM_sub_bytes_0_t32;
reg [4-1:0] FSM_sub_bytes_0_t33;
reg [64-1:0] FSM_sub_bytes_0_t34;
reg [8-1:0] FSM_sub_bytes_0_t35;
reg [64-1:0] FSM_sub_bytes_0_t36;
reg [1024-1:0] FSM_sub_bytes_0_t37;
reg [64-1:0] FSM_sub_bytes_0_t38;
reg [4-1:0] FSM_sub_bytes_0_t39;
reg [64-1:0] FSM_sub_bytes_0_t40;
reg [4-1:0] FSM_sub_bytes_0_t41;
reg [64-1:0] FSM_sub_bytes_0_t42;
reg [8-1:0] FSM_sub_bytes_0_t43;
reg [64-1:0] FSM_sub_bytes_0_t44;
reg [1024-1:0] FSM_sub_bytes_0_t45;
reg [64-1:0] FSM_sub_bytes_0_t46;
reg [4-1:0] FSM_sub_bytes_0_t47;
reg [64-1:0] FSM_sub_bytes_0_t48;
reg [4-1:0] FSM_sub_bytes_0_t49;
reg [64-1:0] FSM_sub_bytes_0_t50;
reg [8-1:0] FSM_sub_bytes_0_t51;
reg [64-1:0] FSM_sub_bytes_0_t52;
reg [1024-1:0] FSM_sub_bytes_0_t53;
reg [64-1:0] FSM_sub_bytes_0_t54;
reg [4-1:0] FSM_sub_bytes_0_t55;
reg [64-1:0] FSM_sub_bytes_0_t56;
reg [4-1:0] FSM_sub_bytes_0_t57;
reg [64-1:0] FSM_sub_bytes_0_t58;
reg [8-1:0] FSM_sub_bytes_0_t59;
reg [64-1:0] FSM_sub_bytes_0_t60;
reg [1024-1:0] FSM_sub_bytes_0_t61;
reg [64-1:0] FSM_sub_bytes_0_t62;
reg [4-1:0] FSM_sub_bytes_0_t63;
reg [64-1:0] FSM_sub_bytes_0_t64;
reg [4-1:0] FSM_sub_bytes_0_t65;
reg [64-1:0] FSM_sub_bytes_0_t66;
reg [8-1:0] FSM_sub_bytes_0_t67;
reg [64-1:0] FSM_sub_bytes_0_t68;
reg [1024-1:0] FSM_sub_bytes_0_t69;
reg [64-1:0] FSM_sub_bytes_0_t70;
reg [4-1:0] FSM_sub_bytes_0_t71;
reg [64-1:0] FSM_sub_bytes_0_t72;
reg [4-1:0] FSM_sub_bytes_0_t73;
reg [64-1:0] FSM_sub_bytes_0_t74;
reg [8-1:0] FSM_sub_bytes_0_t75;
reg [64-1:0] FSM_sub_bytes_0_t76;
reg [1024-1:0] FSM_sub_bytes_0_t77;
reg [64-1:0] FSM_sub_bytes_0_t78;
reg [4-1:0] FSM_sub_bytes_0_t79;
reg [64-1:0] FSM_sub_bytes_0_t80;
reg [4-1:0] FSM_sub_bytes_0_t81;
reg [64-1:0] FSM_sub_bytes_0_t82;
reg [8-1:0] FSM_sub_bytes_0_t83;
reg [64-1:0] FSM_sub_bytes_0_t84;
reg [1024-1:0] FSM_sub_bytes_0_t85;
reg [64-1:0] FSM_sub_bytes_0_t86;
reg [4-1:0] FSM_sub_bytes_0_t87;
reg [64-1:0] FSM_sub_bytes_0_t88;
reg [4-1:0] FSM_sub_bytes_0_t89;
reg [64-1:0] FSM_sub_bytes_0_t90;
reg [8-1:0] FSM_sub_bytes_0_t91;
reg [64-1:0] FSM_sub_bytes_0_t92;
reg [1024-1:0] FSM_sub_bytes_0_t93;
reg [64-1:0] FSM_sub_bytes_0_t94;
reg [4-1:0] FSM_sub_bytes_0_t95;
reg [64-1:0] FSM_sub_bytes_0_t96;
reg [4-1:0] FSM_sub_bytes_0_t97;
reg [64-1:0] FSM_sub_bytes_0_t98;
reg [8-1:0] FSM_sub_bytes_0_t99;
reg [64-1:0] FSM_sub_bytes_0_t100;
reg [1024-1:0] FSM_sub_bytes_0_t101;
reg [64-1:0] FSM_sub_bytes_0_t102;
reg [4-1:0] FSM_sub_bytes_0_t103;
reg [64-1:0] FSM_sub_bytes_0_t104;
reg [4-1:0] FSM_sub_bytes_0_t105;
reg [64-1:0] FSM_sub_bytes_0_t106;
reg [8-1:0] FSM_sub_bytes_0_t107;
reg [64-1:0] FSM_sub_bytes_0_t108;
reg [1024-1:0] FSM_sub_bytes_0_t109;
reg [64-1:0] FSM_sub_bytes_0_t110;
reg [4-1:0] FSM_sub_bytes_0_t111;
reg [64-1:0] FSM_sub_bytes_0_t112;
reg [4-1:0] FSM_sub_bytes_0_t113;
reg [64-1:0] FSM_sub_bytes_0_t114;
reg [8-1:0] FSM_sub_bytes_0_t115;
reg [64-1:0] FSM_sub_bytes_0_t116;
reg [1024-1:0] FSM_sub_bytes_0_t117;
reg [64-1:0] FSM_sub_bytes_0_t118;
reg [4-1:0] FSM_sub_bytes_0_t119;
reg [64-1:0] FSM_sub_bytes_0_t120;
reg [4-1:0] FSM_sub_bytes_0_t121;
reg [64-1:0] FSM_sub_bytes_0_t122;
reg [8-1:0] FSM_sub_bytes_0_t123;
reg [64-1:0] FSM_sub_bytes_0_t124;
reg [1024-1:0] FSM_sub_bytes_0_t125;
reg [64-1:0] FSM_sub_bytes_0_t126;
reg [4-1:0] FSM_sub_bytes_0_t127;
reg [64-1:0] FSM_sub_bytes_0_t128;
reg [4-1:0] FSM_sub_bytes_0_t129;
reg [64-1:0] FSM_sub_bytes_0_t130;
reg [8-1:0] FSM_sub_bytes_0_t131;
reg [64-1:0] FSM_sub_bytes_0_t132;
reg [1024-1:0] FSM_sub_bytes_0_t133;
reg [64-1:0] FSM_sub_bytes_0_t134;
reg [4-1:0] FSM_sub_bytes_0_t135;
reg [64-1:0] FSM_sub_bytes_0_t136;
reg [4-1:0] FSM_sub_bytes_0_t137;
reg [64-1:0] FSM_sub_bytes_0_t138;
reg [8-1:0] FSM_sub_bytes_0_t139;
reg [64-1:0] FSM_sub_bytes_0_t140;
reg [1024-1:0] FSM_sub_bytes_0_t141;
reg [64-1:0] FSM_sub_bytes_0_t142;
reg [4-1:0] FSM_sub_bytes_0_t143;
reg [64-1:0] FSM_sub_bytes_0_t144;
reg [4-1:0] FSM_sub_bytes_0_t145;
reg [64-1:0] FSM_sub_bytes_0_t146;
reg [8-1:0] FSM_sub_bytes_0_t147;
reg [64-1:0] FSM_sub_bytes_0_t148;
reg [1024-1:0] FSM_sub_bytes_0_t149;
reg [64-1:0] FSM_sub_bytes_0_t150;
reg [4-1:0] FSM_sub_bytes_0_t151;
reg [64-1:0] FSM_sub_bytes_0_t152;
reg [4-1:0] FSM_sub_bytes_0_t153;
reg [64-1:0] FSM_sub_bytes_0_t154;
reg [8-1:0] FSM_sub_bytes_0_t155;
reg [64-1:0] FSM_sub_bytes_0_t156;
reg [1024-1:0] FSM_sub_bytes_0_t157;
reg [64-1:0] FSM_sub_bytes_0_t158;
reg [4-1:0] FSM_sub_bytes_0_t159;
reg [64-1:0] FSM_sub_bytes_0_t160;
reg [64-1:0] FSM_sub_bytes_0_t161;
reg [4-1:0] FSM_sub_bytes_0_t162;
reg [64-1:0] FSM_sub_bytes_0_t163;
reg [64-1:0] FSM_sub_bytes_0_t164;
reg [6-1:0] FSM_sub_bytes_0_t165;
reg [64-1:0] FSM_sub_bytes_0_t166;
reg [4-1:0] FSM_sub_bytes_0_t167;
reg [64-1:0] FSM_sub_bytes_0_t168;
reg [64-1:0] FSM_sub_bytes_0_t169;
reg [6-1:0] FSM_sub_bytes_0_t170;
reg [64-1:0] FSM_sub_bytes_0_t171;
reg [4-1:0] FSM_sub_bytes_0_t172;
reg [64-1:0] FSM_sub_bytes_0_t173;
reg [64-1:0] FSM_sub_bytes_0_t174;
reg [6-1:0] FSM_sub_bytes_0_t175;
reg [64-1:0] FSM_sub_bytes_0_t176;
reg [4-1:0] FSM_sub_bytes_0_t177;
reg [64-1:0] FSM_sub_bytes_0_t178;
reg [64-1:0] FSM_sub_bytes_0_t179;
reg [6-1:0] FSM_sub_bytes_0_t180;
reg [64-1:0] FSM_sub_bytes_0_t181;
reg [4-1:0] FSM_sub_bytes_0_t182;
reg [64-1:0] FSM_sub_bytes_0_t183;
reg [64-1:0] FSM_sub_bytes_0_t184;
reg [6-1:0] FSM_sub_bytes_0_t185;
reg [64-1:0] FSM_sub_bytes_0_t186;
reg [4-1:0] FSM_sub_bytes_0_t187;
reg [64-1:0] FSM_sub_bytes_0_t188;
reg [64-1:0] FSM_sub_bytes_0_t189;
reg [6-1:0] FSM_sub_bytes_0_t190;
reg [64-1:0] FSM_sub_bytes_0_t191;
reg [4-1:0] FSM_sub_bytes_0_t192;
reg [64-1:0] FSM_sub_bytes_0_t193;
reg [64-1:0] FSM_sub_bytes_0_t194;
reg [6-1:0] FSM_sub_bytes_0_t195;
reg [64-1:0] FSM_sub_bytes_0_t196;
reg [4-1:0] FSM_sub_bytes_0_t197;
reg [64-1:0] FSM_sub_bytes_0_t198;
reg [64-1:0] FSM_sub_bytes_0_t199;
reg [4-1:0] FSM_sub_bytes_0_t200;
reg [64-1:0] FSM_sub_bytes_0_t201;
reg [64-1:0] FSM_sub_bytes_0_t202;
reg [6-1:0] FSM_sub_bytes_0_t203;
reg [64-1:0] FSM_sub_bytes_0_t204;
reg [4-1:0] FSM_sub_bytes_0_t205;
reg [64-1:0] FSM_sub_bytes_0_t206;
reg [64-1:0] FSM_sub_bytes_0_t207;
reg [6-1:0] FSM_sub_bytes_0_t208;
reg [64-1:0] FSM_sub_bytes_0_t209;
reg [4-1:0] FSM_sub_bytes_0_t210;
reg [64-1:0] FSM_sub_bytes_0_t211;
reg [64-1:0] FSM_sub_bytes_0_t212;
reg [6-1:0] FSM_sub_bytes_0_t213;
reg [64-1:0] FSM_sub_bytes_0_t214;
reg [4-1:0] FSM_sub_bytes_0_t215;
reg [64-1:0] FSM_sub_bytes_0_t216;
reg [64-1:0] FSM_sub_bytes_0_t217;
reg [6-1:0] FSM_sub_bytes_0_t218;
reg [64-1:0] FSM_sub_bytes_0_t219;
reg [4-1:0] FSM_sub_bytes_0_t220;
reg [64-1:0] FSM_sub_bytes_0_t221;
reg [64-1:0] FSM_sub_bytes_0_t222;
reg [6-1:0] FSM_sub_bytes_0_t223;
reg [64-1:0] FSM_sub_bytes_0_t224;
reg [4-1:0] FSM_sub_bytes_0_t225;
reg [64-1:0] FSM_sub_bytes_0_t226;
reg [64-1:0] FSM_sub_bytes_0_t227;
reg [6-1:0] FSM_sub_bytes_0_t228;
reg [64-1:0] FSM_sub_bytes_0_t229;
reg [4-1:0] FSM_sub_bytes_0_t230;
reg [64-1:0] FSM_sub_bytes_0_t231;
reg [64-1:0] FSM_sub_bytes_0_t232;
reg [6-1:0] FSM_sub_bytes_0_t233;

assign FSM_sub_bytes_0_out_higher_out = ((((((FSM_sub_bytes_0_t160 | (FSM_sub_bytes_0_t163 << FSM_sub_bytes_0_t165)) | (FSM_sub_bytes_0_t168 << FSM_sub_bytes_0_t170)) | (FSM_sub_bytes_0_t173 << FSM_sub_bytes_0_t175)) | (FSM_sub_bytes_0_t178 << FSM_sub_bytes_0_t180)) | (FSM_sub_bytes_0_t183 << FSM_sub_bytes_0_t185)) | (FSM_sub_bytes_0_t188 << FSM_sub_bytes_0_t190)) | (FSM_sub_bytes_0_t193 << FSM_sub_bytes_0_t195);
assign FSM_sub_bytes_0_out_lower_out = ((((((FSM_sub_bytes_0_t198 | (FSM_sub_bytes_0_t201 << FSM_sub_bytes_0_t203)) | (FSM_sub_bytes_0_t206 << FSM_sub_bytes_0_t208)) | (FSM_sub_bytes_0_t211 << FSM_sub_bytes_0_t213)) | (FSM_sub_bytes_0_t216 << FSM_sub_bytes_0_t218)) | (FSM_sub_bytes_0_t221 << FSM_sub_bytes_0_t223)) | (FSM_sub_bytes_0_t226 << FSM_sub_bytes_0_t228)) | (FSM_sub_bytes_0_t231 << FSM_sub_bytes_0_t233);
assign FSM_sub_bytes_0_out_valid = 1'b1;


/*
    Wiring by sub_bytes
*/
assign i_ready = FSM_sub_bytes_0_in_ready;
assign o_higher_out = FSM_sub_bytes_0_out_higher_out;
assign o_lower_out = FSM_sub_bytes_0_out_lower_out;
assign o_valid = FSM_sub_bytes_0_out_valid;
/* End wiring by sub_bytes */


initial begin
    FSM_sub_bytes_0_t0[0 * 64 +: 64] = i_lower_bits & 64'b0000000000000000000000000000000000000000000000000000000011111111;
    FSM_sub_bytes_0_t1 = 64'b0000000000000000000000000000000000000000000000000000000000001000;
    FSM_sub_bytes_0_t2 = FSM_sub_bytes_0_t1[6'b0 * 1 +: 6 * 1];
    FSM_sub_bytes_0_t0[1 * 64 +: 64] = (i_lower_bits >> FSM_sub_bytes_0_t2) & 64'b0000000000000000000000000000000000000000000000000000000011111111;
    FSM_sub_bytes_0_t3 = 64'b0000000000000000000000000000000000000000000000000000000000010000;
    FSM_sub_bytes_0_t4 = FSM_sub_bytes_0_t3[6'b0 * 1 +: 6 * 1];
    FSM_sub_bytes_0_t0[2 * 64 +: 64] = (i_lower_bits >> FSM_sub_bytes_0_t4) & 64'b0000000000000000000000000000000000000000000000000000000011111111;
    FSM_sub_bytes_0_t5 = 64'b0000000000000000000000000000000000000000000000000000000000011000;
    FSM_sub_bytes_0_t6 = FSM_sub_bytes_0_t5[6'b0 * 1 +: 6 * 1];
    FSM_sub_bytes_0_t0[3 * 64 +: 64] = (i_lower_bits >> FSM_sub_bytes_0_t6) & 64'b0000000000000000000000000000000000000000000000000000000011111111;
    FSM_sub_bytes_0_t7 = 64'b0000000000000000000000000000000000000000000000000000000000100000;
    FSM_sub_bytes_0_t8 = FSM_sub_bytes_0_t7[6'b0 * 1 +: 6 * 1];
    FSM_sub_bytes_0_t0[4 * 64 +: 64] = (i_lower_bits >> FSM_sub_bytes_0_t8) & 64'b0000000000000000000000000000000000000000000000000000000011111111;
    FSM_sub_bytes_0_t9 = 64'b0000000000000000000000000000000000000000000000000000000000101000;
    FSM_sub_bytes_0_t10 = FSM_sub_bytes_0_t9[6'b0 * 1 +: 6 * 1];
    FSM_sub_bytes_0_t0[5 * 64 +: 64] = (i_lower_bits >> FSM_sub_bytes_0_t10) & 64'b0000000000000000000000000000000000000000000000000000000011111111;
    FSM_sub_bytes_0_t11 = 64'b0000000000000000000000000000000000000000000000000000000000110000;
    FSM_sub_bytes_0_t12 = FSM_sub_bytes_0_t11[6'b0 * 1 +: 6 * 1];
    FSM_sub_bytes_0_t0[6 * 64 +: 64] = (i_lower_bits >> FSM_sub_bytes_0_t12) & 64'b0000000000000000000000000000000000000000000000000000000011111111;
    FSM_sub_bytes_0_t13 = 64'b0000000000000000000000000000000000000000000000000000000000111000;
    FSM_sub_bytes_0_t14 = FSM_sub_bytes_0_t13[6'b0 * 1 +: 6 * 1];
    FSM_sub_bytes_0_t0[7 * 64 +: 64] = (i_lower_bits >> FSM_sub_bytes_0_t14) & 64'b0000000000000000000000000000000000000000000000000000000011111111;
    FSM_sub_bytes_0_t0[8 * 64 +: 64] = i_higher_bits & 64'b0000000000000000000000000000000000000000000000000000000011111111;
    FSM_sub_bytes_0_t15 = 64'b0000000000000000000000000000000000000000000000000000000000001000;
    FSM_sub_bytes_0_t16 = FSM_sub_bytes_0_t15[6'b0 * 1 +: 6 * 1];
    FSM_sub_bytes_0_t0[9 * 64 +: 64] = (i_higher_bits >> FSM_sub_bytes_0_t16) & 64'b0000000000000000000000000000000000000000000000000000000011111111;
    FSM_sub_bytes_0_t17 = 64'b0000000000000000000000000000000000000000000000000000000000010000;
    FSM_sub_bytes_0_t18 = FSM_sub_bytes_0_t17[6'b0 * 1 +: 6 * 1];
    FSM_sub_bytes_0_t0[10 * 64 +: 64] = (i_higher_bits >> FSM_sub_bytes_0_t18) & 64'b0000000000000000000000000000000000000000000000000000000011111111;
    FSM_sub_bytes_0_t19 = 64'b0000000000000000000000000000000000000000000000000000000000011000;
    FSM_sub_bytes_0_t20 = FSM_sub_bytes_0_t19[6'b0 * 1 +: 6 * 1];
    FSM_sub_bytes_0_t0[11 * 64 +: 64] = (i_higher_bits >> FSM_sub_bytes_0_t20) & 64'b0000000000000000000000000000000000000000000000000000000011111111;
    FSM_sub_bytes_0_t21 = 64'b0000000000000000000000000000000000000000000000000000000000100000;
    FSM_sub_bytes_0_t22 = FSM_sub_bytes_0_t21[6'b0 * 1 +: 6 * 1];
    FSM_sub_bytes_0_t0[12 * 64 +: 64] = (i_higher_bits >> FSM_sub_bytes_0_t22) & 64'b0000000000000000000000000000000000000000000000000000000011111111;
    FSM_sub_bytes_0_t23 = 64'b0000000000000000000000000000000000000000000000000000000000101000;
    FSM_sub_bytes_0_t24 = FSM_sub_bytes_0_t23[6'b0 * 1 +: 6 * 1];
    FSM_sub_bytes_0_t0[13 * 64 +: 64] = (i_higher_bits >> FSM_sub_bytes_0_t24) & 64'b0000000000000000000000000000000000000000000000000000000011111111;
    FSM_sub_bytes_0_t25 = 64'b0000000000000000000000000000000000000000000000000000000000110000;
    FSM_sub_bytes_0_t26 = FSM_sub_bytes_0_t25[6'b0 * 1 +: 6 * 1];
    FSM_sub_bytes_0_t0[14 * 64 +: 64] = (i_higher_bits >> FSM_sub_bytes_0_t26) & 64'b0000000000000000000000000000000000000000000000000000000011111111;
    FSM_sub_bytes_0_t27 = 64'b0000000000000000000000000000000000000000000000000000000000111000;
    FSM_sub_bytes_0_t28 = FSM_sub_bytes_0_t27[6'b0 * 1 +: 6 * 1];
    FSM_sub_bytes_0_t0[15 * 64 +: 64] = (i_higher_bits >> FSM_sub_bytes_0_t28) & 64'b0000000000000000000000000000000000000000000000000000000011111111;
    FSM_sub_bytes_0_t29 = 64'b0;
    FSM_sub_bytes_0_t30 = FSM_sub_bytes_0_t29[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t31[0 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001100011;
    FSM_sub_bytes_0_t31[1 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001111100;
    FSM_sub_bytes_0_t31[2 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001110111;
    FSM_sub_bytes_0_t31[3 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001111011;
    FSM_sub_bytes_0_t31[4 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011110010;
    FSM_sub_bytes_0_t31[5 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001101011;
    FSM_sub_bytes_0_t31[6 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001101111;
    FSM_sub_bytes_0_t31[7 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011000101;
    FSM_sub_bytes_0_t31[8 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000110000;
    FSM_sub_bytes_0_t31[9 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000000001;
    FSM_sub_bytes_0_t31[10 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001100111;
    FSM_sub_bytes_0_t31[11 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000101011;
    FSM_sub_bytes_0_t31[12 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011111110;
    FSM_sub_bytes_0_t31[13 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011010111;
    FSM_sub_bytes_0_t31[14 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010101011;
    FSM_sub_bytes_0_t31[15 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001110110;
    FSM_sub_bytes_0_t31[16 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011001010;
    FSM_sub_bytes_0_t31[17 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010000010;
    FSM_sub_bytes_0_t31[18 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011001001;
    FSM_sub_bytes_0_t31[19 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001111101;
    FSM_sub_bytes_0_t31[20 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011111010;
    FSM_sub_bytes_0_t31[21 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001011001;
    FSM_sub_bytes_0_t31[22 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001000111;
    FSM_sub_bytes_0_t31[23 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011110000;
    FSM_sub_bytes_0_t31[24 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010101101;
    FSM_sub_bytes_0_t31[25 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011010100;
    FSM_sub_bytes_0_t31[26 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010100010;
    FSM_sub_bytes_0_t31[27 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010101111;
    FSM_sub_bytes_0_t31[28 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010011100;
    FSM_sub_bytes_0_t31[29 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010100100;
    FSM_sub_bytes_0_t31[30 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001110010;
    FSM_sub_bytes_0_t31[31 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011000000;
    FSM_sub_bytes_0_t31[32 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010110111;
    FSM_sub_bytes_0_t31[33 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011111101;
    FSM_sub_bytes_0_t31[34 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010010011;
    FSM_sub_bytes_0_t31[35 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000100110;
    FSM_sub_bytes_0_t31[36 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000110110;
    FSM_sub_bytes_0_t31[37 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000111111;
    FSM_sub_bytes_0_t31[38 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011110111;
    FSM_sub_bytes_0_t31[39 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011001100;
    FSM_sub_bytes_0_t31[40 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000110100;
    FSM_sub_bytes_0_t31[41 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010100101;
    FSM_sub_bytes_0_t31[42 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011100101;
    FSM_sub_bytes_0_t31[43 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011110001;
    FSM_sub_bytes_0_t31[44 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001110001;
    FSM_sub_bytes_0_t31[45 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011011000;
    FSM_sub_bytes_0_t31[46 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000110001;
    FSM_sub_bytes_0_t31[47 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000010101;
    FSM_sub_bytes_0_t31[48 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000000100;
    FSM_sub_bytes_0_t31[49 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011000111;
    FSM_sub_bytes_0_t31[50 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000100011;
    FSM_sub_bytes_0_t31[51 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011000011;
    FSM_sub_bytes_0_t31[52 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000011000;
    FSM_sub_bytes_0_t31[53 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010010110;
    FSM_sub_bytes_0_t31[54 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000000101;
    FSM_sub_bytes_0_t31[55 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010011010;
    FSM_sub_bytes_0_t31[56 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000000111;
    FSM_sub_bytes_0_t31[57 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000010010;
    FSM_sub_bytes_0_t31[58 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010000000;
    FSM_sub_bytes_0_t31[59 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011100010;
    FSM_sub_bytes_0_t31[60 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011101011;
    FSM_sub_bytes_0_t31[61 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000100111;
    FSM_sub_bytes_0_t31[62 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010110010;
    FSM_sub_bytes_0_t31[63 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001110101;
    FSM_sub_bytes_0_t31[64 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000001001;
    FSM_sub_bytes_0_t31[65 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010000011;
    FSM_sub_bytes_0_t31[66 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000101100;
    FSM_sub_bytes_0_t31[67 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000011010;
    FSM_sub_bytes_0_t31[68 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000011011;
    FSM_sub_bytes_0_t31[69 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001101110;
    FSM_sub_bytes_0_t31[70 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001011010;
    FSM_sub_bytes_0_t31[71 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010100000;
    FSM_sub_bytes_0_t31[72 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001010010;
    FSM_sub_bytes_0_t31[73 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000111011;
    FSM_sub_bytes_0_t31[74 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011010110;
    FSM_sub_bytes_0_t31[75 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010110011;
    FSM_sub_bytes_0_t31[76 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000101001;
    FSM_sub_bytes_0_t31[77 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011100011;
    FSM_sub_bytes_0_t31[78 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000101111;
    FSM_sub_bytes_0_t31[79 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010000100;
    FSM_sub_bytes_0_t31[80 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001010011;
    FSM_sub_bytes_0_t31[81 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011010001;
    FSM_sub_bytes_0_t31[82 * 64 +: 64] = 64'b0;
    FSM_sub_bytes_0_t31[83 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011101101;
    FSM_sub_bytes_0_t31[84 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000100000;
    FSM_sub_bytes_0_t31[85 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011111100;
    FSM_sub_bytes_0_t31[86 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010110001;
    FSM_sub_bytes_0_t31[87 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001011011;
    FSM_sub_bytes_0_t31[88 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001101010;
    FSM_sub_bytes_0_t31[89 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011001011;
    FSM_sub_bytes_0_t31[90 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010111110;
    FSM_sub_bytes_0_t31[91 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000111001;
    FSM_sub_bytes_0_t31[92 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001001010;
    FSM_sub_bytes_0_t31[93 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001001100;
    FSM_sub_bytes_0_t31[94 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001011000;
    FSM_sub_bytes_0_t31[95 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011001111;
    FSM_sub_bytes_0_t31[96 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011010000;
    FSM_sub_bytes_0_t31[97 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011101111;
    FSM_sub_bytes_0_t31[98 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010101010;
    FSM_sub_bytes_0_t31[99 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011111011;
    FSM_sub_bytes_0_t31[100 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001000011;
    FSM_sub_bytes_0_t31[101 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001001101;
    FSM_sub_bytes_0_t31[102 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000110011;
    FSM_sub_bytes_0_t31[103 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010000101;
    FSM_sub_bytes_0_t31[104 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001000101;
    FSM_sub_bytes_0_t31[105 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011111001;
    FSM_sub_bytes_0_t31[106 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000000010;
    FSM_sub_bytes_0_t31[107 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001111111;
    FSM_sub_bytes_0_t31[108 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001010000;
    FSM_sub_bytes_0_t31[109 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000111100;
    FSM_sub_bytes_0_t31[110 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010011111;
    FSM_sub_bytes_0_t31[111 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010101000;
    FSM_sub_bytes_0_t31[112 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001010001;
    FSM_sub_bytes_0_t31[113 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010100011;
    FSM_sub_bytes_0_t31[114 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001000000;
    FSM_sub_bytes_0_t31[115 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010001111;
    FSM_sub_bytes_0_t31[116 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010010010;
    FSM_sub_bytes_0_t31[117 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010011101;
    FSM_sub_bytes_0_t31[118 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000111000;
    FSM_sub_bytes_0_t31[119 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011110101;
    FSM_sub_bytes_0_t31[120 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010111100;
    FSM_sub_bytes_0_t31[121 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010110110;
    FSM_sub_bytes_0_t31[122 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011011010;
    FSM_sub_bytes_0_t31[123 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000100001;
    FSM_sub_bytes_0_t31[124 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000010000;
    FSM_sub_bytes_0_t31[125 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011111111;
    FSM_sub_bytes_0_t31[126 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011110011;
    FSM_sub_bytes_0_t31[127 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011010010;
    FSM_sub_bytes_0_t31[128 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011001101;
    FSM_sub_bytes_0_t31[129 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000001100;
    FSM_sub_bytes_0_t31[130 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000010011;
    FSM_sub_bytes_0_t31[131 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011101100;
    FSM_sub_bytes_0_t31[132 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001011111;
    FSM_sub_bytes_0_t31[133 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010010111;
    FSM_sub_bytes_0_t31[134 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001000100;
    FSM_sub_bytes_0_t31[135 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000010111;
    FSM_sub_bytes_0_t31[136 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011000100;
    FSM_sub_bytes_0_t31[137 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010100111;
    FSM_sub_bytes_0_t31[138 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001111110;
    FSM_sub_bytes_0_t31[139 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000111101;
    FSM_sub_bytes_0_t31[140 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001100100;
    FSM_sub_bytes_0_t31[141 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001011101;
    FSM_sub_bytes_0_t31[142 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000011001;
    FSM_sub_bytes_0_t31[143 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001110011;
    FSM_sub_bytes_0_t31[144 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001100000;
    FSM_sub_bytes_0_t31[145 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010000001;
    FSM_sub_bytes_0_t31[146 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001001111;
    FSM_sub_bytes_0_t31[147 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011011100;
    FSM_sub_bytes_0_t31[148 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000100010;
    FSM_sub_bytes_0_t31[149 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000101010;
    FSM_sub_bytes_0_t31[150 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010010000;
    FSM_sub_bytes_0_t31[151 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010001000;
    FSM_sub_bytes_0_t31[152 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001000110;
    FSM_sub_bytes_0_t31[153 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011101110;
    FSM_sub_bytes_0_t31[154 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010111000;
    FSM_sub_bytes_0_t31[155 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000010100;
    FSM_sub_bytes_0_t31[156 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011011110;
    FSM_sub_bytes_0_t31[157 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001011110;
    FSM_sub_bytes_0_t31[158 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000001011;
    FSM_sub_bytes_0_t31[159 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011011011;
    FSM_sub_bytes_0_t31[160 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011100000;
    FSM_sub_bytes_0_t31[161 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000110010;
    FSM_sub_bytes_0_t31[162 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000111010;
    FSM_sub_bytes_0_t31[163 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000001010;
    FSM_sub_bytes_0_t31[164 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001001001;
    FSM_sub_bytes_0_t31[165 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000000110;
    FSM_sub_bytes_0_t31[166 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000100100;
    FSM_sub_bytes_0_t31[167 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001011100;
    FSM_sub_bytes_0_t31[168 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011000010;
    FSM_sub_bytes_0_t31[169 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011010011;
    FSM_sub_bytes_0_t31[170 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010101100;
    FSM_sub_bytes_0_t31[171 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001100010;
    FSM_sub_bytes_0_t31[172 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010010001;
    FSM_sub_bytes_0_t31[173 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010010101;
    FSM_sub_bytes_0_t31[174 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011100100;
    FSM_sub_bytes_0_t31[175 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001111001;
    FSM_sub_bytes_0_t31[176 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011100111;
    FSM_sub_bytes_0_t31[177 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011001000;
    FSM_sub_bytes_0_t31[178 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000110111;
    FSM_sub_bytes_0_t31[179 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001101101;
    FSM_sub_bytes_0_t31[180 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010001101;
    FSM_sub_bytes_0_t31[181 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011010101;
    FSM_sub_bytes_0_t31[182 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001001110;
    FSM_sub_bytes_0_t31[183 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010101001;
    FSM_sub_bytes_0_t31[184 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001101100;
    FSM_sub_bytes_0_t31[185 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001010110;
    FSM_sub_bytes_0_t31[186 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011110100;
    FSM_sub_bytes_0_t31[187 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011101010;
    FSM_sub_bytes_0_t31[188 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001100101;
    FSM_sub_bytes_0_t31[189 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001111010;
    FSM_sub_bytes_0_t31[190 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010101110;
    FSM_sub_bytes_0_t31[191 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000001000;
    FSM_sub_bytes_0_t31[192 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010111010;
    FSM_sub_bytes_0_t31[193 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001111000;
    FSM_sub_bytes_0_t31[194 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000100101;
    FSM_sub_bytes_0_t31[195 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000101110;
    FSM_sub_bytes_0_t31[196 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000011100;
    FSM_sub_bytes_0_t31[197 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010100110;
    FSM_sub_bytes_0_t31[198 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010110100;
    FSM_sub_bytes_0_t31[199 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011000110;
    FSM_sub_bytes_0_t31[200 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011101000;
    FSM_sub_bytes_0_t31[201 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011011101;
    FSM_sub_bytes_0_t31[202 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001110100;
    FSM_sub_bytes_0_t31[203 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000011111;
    FSM_sub_bytes_0_t31[204 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001001011;
    FSM_sub_bytes_0_t31[205 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010111101;
    FSM_sub_bytes_0_t31[206 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010001011;
    FSM_sub_bytes_0_t31[207 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010001010;
    FSM_sub_bytes_0_t31[208 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001110000;
    FSM_sub_bytes_0_t31[209 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000111110;
    FSM_sub_bytes_0_t31[210 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010110101;
    FSM_sub_bytes_0_t31[211 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001100110;
    FSM_sub_bytes_0_t31[212 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001001000;
    FSM_sub_bytes_0_t31[213 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000000011;
    FSM_sub_bytes_0_t31[214 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011110110;
    FSM_sub_bytes_0_t31[215 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000001110;
    FSM_sub_bytes_0_t31[216 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001100001;
    FSM_sub_bytes_0_t31[217 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000110101;
    FSM_sub_bytes_0_t31[218 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001010111;
    FSM_sub_bytes_0_t31[219 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010111001;
    FSM_sub_bytes_0_t31[220 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010000110;
    FSM_sub_bytes_0_t31[221 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011000001;
    FSM_sub_bytes_0_t31[222 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000011101;
    FSM_sub_bytes_0_t31[223 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010011110;
    FSM_sub_bytes_0_t31[224 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011100001;
    FSM_sub_bytes_0_t31[225 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011111000;
    FSM_sub_bytes_0_t31[226 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010011000;
    FSM_sub_bytes_0_t31[227 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000010001;
    FSM_sub_bytes_0_t31[228 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001101001;
    FSM_sub_bytes_0_t31[229 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011011001;
    FSM_sub_bytes_0_t31[230 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010001110;
    FSM_sub_bytes_0_t31[231 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010010100;
    FSM_sub_bytes_0_t31[232 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010011011;
    FSM_sub_bytes_0_t31[233 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000011110;
    FSM_sub_bytes_0_t31[234 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010000111;
    FSM_sub_bytes_0_t31[235 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011101001;
    FSM_sub_bytes_0_t31[236 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011001110;
    FSM_sub_bytes_0_t31[237 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001010101;
    FSM_sub_bytes_0_t31[238 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000101000;
    FSM_sub_bytes_0_t31[239 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011011111;
    FSM_sub_bytes_0_t31[240 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010001100;
    FSM_sub_bytes_0_t31[241 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010100001;
    FSM_sub_bytes_0_t31[242 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010001001;
    FSM_sub_bytes_0_t31[243 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000001101;
    FSM_sub_bytes_0_t31[244 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010111111;
    FSM_sub_bytes_0_t31[245 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011100110;
    FSM_sub_bytes_0_t31[246 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001000010;
    FSM_sub_bytes_0_t31[247 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001101000;
    FSM_sub_bytes_0_t31[248 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001000001;
    FSM_sub_bytes_0_t31[249 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010011001;
    FSM_sub_bytes_0_t31[250 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000101101;
    FSM_sub_bytes_0_t31[251 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000001111;
    FSM_sub_bytes_0_t31[252 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010110000;
    FSM_sub_bytes_0_t31[253 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001010100;
    FSM_sub_bytes_0_t31[254 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010111011;
    FSM_sub_bytes_0_t31[255 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000010110;
    FSM_sub_bytes_0_t32 = 64'b0;
    FSM_sub_bytes_0_t33 = FSM_sub_bytes_0_t32[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t34 = FSM_sub_bytes_0_t0[FSM_sub_bytes_0_t33 * 64 +: 64];
    FSM_sub_bytes_0_t35 = FSM_sub_bytes_0_t34[6'b0 * 1 +: 8 * 1];
    FSM_sub_bytes_0_t36 = FSM_sub_bytes_0_t31[FSM_sub_bytes_0_t35 * 64 +: 64];
    FSM_sub_bytes_0_t37 = FSM_sub_bytes_0_t0;
    FSM_sub_bytes_0_t37[FSM_sub_bytes_0_t30 * 64 +: 64] = FSM_sub_bytes_0_t36;
    FSM_sub_bytes_0_t38 = 64'b0000000000000000000000000000000000000000000000000000000000000001;
    FSM_sub_bytes_0_t39 = FSM_sub_bytes_0_t38[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t40 = 64'b0000000000000000000000000000000000000000000000000000000000000001;
    FSM_sub_bytes_0_t41 = FSM_sub_bytes_0_t40[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t42 = FSM_sub_bytes_0_t37[FSM_sub_bytes_0_t41 * 64 +: 64];
    FSM_sub_bytes_0_t43 = FSM_sub_bytes_0_t42[6'b0 * 1 +: 8 * 1];
    FSM_sub_bytes_0_t44 = FSM_sub_bytes_0_t31[FSM_sub_bytes_0_t43 * 64 +: 64];
    FSM_sub_bytes_0_t45 = FSM_sub_bytes_0_t37;
    FSM_sub_bytes_0_t45[FSM_sub_bytes_0_t39 * 64 +: 64] = FSM_sub_bytes_0_t44;
    FSM_sub_bytes_0_t46 = 64'b0000000000000000000000000000000000000000000000000000000000000010;
    FSM_sub_bytes_0_t47 = FSM_sub_bytes_0_t46[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t48 = 64'b0000000000000000000000000000000000000000000000000000000000000010;
    FSM_sub_bytes_0_t49 = FSM_sub_bytes_0_t48[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t50 = FSM_sub_bytes_0_t45[FSM_sub_bytes_0_t49 * 64 +: 64];
    FSM_sub_bytes_0_t51 = FSM_sub_bytes_0_t50[6'b0 * 1 +: 8 * 1];
    FSM_sub_bytes_0_t52 = FSM_sub_bytes_0_t31[FSM_sub_bytes_0_t51 * 64 +: 64];
    FSM_sub_bytes_0_t53 = FSM_sub_bytes_0_t45;
    FSM_sub_bytes_0_t53[FSM_sub_bytes_0_t47 * 64 +: 64] = FSM_sub_bytes_0_t52;
    FSM_sub_bytes_0_t54 = 64'b0000000000000000000000000000000000000000000000000000000000000011;
    FSM_sub_bytes_0_t55 = FSM_sub_bytes_0_t54[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t56 = 64'b0000000000000000000000000000000000000000000000000000000000000011;
    FSM_sub_bytes_0_t57 = FSM_sub_bytes_0_t56[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t58 = FSM_sub_bytes_0_t53[FSM_sub_bytes_0_t57 * 64 +: 64];
    FSM_sub_bytes_0_t59 = FSM_sub_bytes_0_t58[6'b0 * 1 +: 8 * 1];
    FSM_sub_bytes_0_t60 = FSM_sub_bytes_0_t31[FSM_sub_bytes_0_t59 * 64 +: 64];
    FSM_sub_bytes_0_t61 = FSM_sub_bytes_0_t53;
    FSM_sub_bytes_0_t61[FSM_sub_bytes_0_t55 * 64 +: 64] = FSM_sub_bytes_0_t60;
    FSM_sub_bytes_0_t62 = 64'b0000000000000000000000000000000000000000000000000000000000000100;
    FSM_sub_bytes_0_t63 = FSM_sub_bytes_0_t62[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t64 = 64'b0000000000000000000000000000000000000000000000000000000000000100;
    FSM_sub_bytes_0_t65 = FSM_sub_bytes_0_t64[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t66 = FSM_sub_bytes_0_t61[FSM_sub_bytes_0_t65 * 64 +: 64];
    FSM_sub_bytes_0_t67 = FSM_sub_bytes_0_t66[6'b0 * 1 +: 8 * 1];
    FSM_sub_bytes_0_t68 = FSM_sub_bytes_0_t31[FSM_sub_bytes_0_t67 * 64 +: 64];
    FSM_sub_bytes_0_t69 = FSM_sub_bytes_0_t61;
    FSM_sub_bytes_0_t69[FSM_sub_bytes_0_t63 * 64 +: 64] = FSM_sub_bytes_0_t68;
    FSM_sub_bytes_0_t70 = 64'b0000000000000000000000000000000000000000000000000000000000000101;
    FSM_sub_bytes_0_t71 = FSM_sub_bytes_0_t70[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t72 = 64'b0000000000000000000000000000000000000000000000000000000000000101;
    FSM_sub_bytes_0_t73 = FSM_sub_bytes_0_t72[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t74 = FSM_sub_bytes_0_t69[FSM_sub_bytes_0_t73 * 64 +: 64];
    FSM_sub_bytes_0_t75 = FSM_sub_bytes_0_t74[6'b0 * 1 +: 8 * 1];
    FSM_sub_bytes_0_t76 = FSM_sub_bytes_0_t31[FSM_sub_bytes_0_t75 * 64 +: 64];
    FSM_sub_bytes_0_t77 = FSM_sub_bytes_0_t69;
    FSM_sub_bytes_0_t77[FSM_sub_bytes_0_t71 * 64 +: 64] = FSM_sub_bytes_0_t76;
    FSM_sub_bytes_0_t78 = 64'b0000000000000000000000000000000000000000000000000000000000000110;
    FSM_sub_bytes_0_t79 = FSM_sub_bytes_0_t78[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t80 = 64'b0000000000000000000000000000000000000000000000000000000000000110;
    FSM_sub_bytes_0_t81 = FSM_sub_bytes_0_t80[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t82 = FSM_sub_bytes_0_t77[FSM_sub_bytes_0_t81 * 64 +: 64];
    FSM_sub_bytes_0_t83 = FSM_sub_bytes_0_t82[6'b0 * 1 +: 8 * 1];
    FSM_sub_bytes_0_t84 = FSM_sub_bytes_0_t31[FSM_sub_bytes_0_t83 * 64 +: 64];
    FSM_sub_bytes_0_t85 = FSM_sub_bytes_0_t77;
    FSM_sub_bytes_0_t85[FSM_sub_bytes_0_t79 * 64 +: 64] = FSM_sub_bytes_0_t84;
    FSM_sub_bytes_0_t86 = 64'b0000000000000000000000000000000000000000000000000000000000000111;
    FSM_sub_bytes_0_t87 = FSM_sub_bytes_0_t86[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t88 = 64'b0000000000000000000000000000000000000000000000000000000000000111;
    FSM_sub_bytes_0_t89 = FSM_sub_bytes_0_t88[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t90 = FSM_sub_bytes_0_t85[FSM_sub_bytes_0_t89 * 64 +: 64];
    FSM_sub_bytes_0_t91 = FSM_sub_bytes_0_t90[6'b0 * 1 +: 8 * 1];
    FSM_sub_bytes_0_t92 = FSM_sub_bytes_0_t31[FSM_sub_bytes_0_t91 * 64 +: 64];
    FSM_sub_bytes_0_t93 = FSM_sub_bytes_0_t85;
    FSM_sub_bytes_0_t93[FSM_sub_bytes_0_t87 * 64 +: 64] = FSM_sub_bytes_0_t92;
    FSM_sub_bytes_0_t94 = 64'b0000000000000000000000000000000000000000000000000000000000001000;
    FSM_sub_bytes_0_t95 = FSM_sub_bytes_0_t94[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t96 = 64'b0000000000000000000000000000000000000000000000000000000000001000;
    FSM_sub_bytes_0_t97 = FSM_sub_bytes_0_t96[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t98 = FSM_sub_bytes_0_t93[FSM_sub_bytes_0_t97 * 64 +: 64];
    FSM_sub_bytes_0_t99 = FSM_sub_bytes_0_t98[6'b0 * 1 +: 8 * 1];
    FSM_sub_bytes_0_t100 = FSM_sub_bytes_0_t31[FSM_sub_bytes_0_t99 * 64 +: 64];
    FSM_sub_bytes_0_t101 = FSM_sub_bytes_0_t93;
    FSM_sub_bytes_0_t101[FSM_sub_bytes_0_t95 * 64 +: 64] = FSM_sub_bytes_0_t100;
    FSM_sub_bytes_0_t102 = 64'b0000000000000000000000000000000000000000000000000000000000001001;
    FSM_sub_bytes_0_t103 = FSM_sub_bytes_0_t102[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t104 = 64'b0000000000000000000000000000000000000000000000000000000000001001;
    FSM_sub_bytes_0_t105 = FSM_sub_bytes_0_t104[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t106 = FSM_sub_bytes_0_t101[FSM_sub_bytes_0_t105 * 64 +: 64];
    FSM_sub_bytes_0_t107 = FSM_sub_bytes_0_t106[6'b0 * 1 +: 8 * 1];
    FSM_sub_bytes_0_t108 = FSM_sub_bytes_0_t31[FSM_sub_bytes_0_t107 * 64 +: 64];
    FSM_sub_bytes_0_t109 = FSM_sub_bytes_0_t101;
    FSM_sub_bytes_0_t109[FSM_sub_bytes_0_t103 * 64 +: 64] = FSM_sub_bytes_0_t108;
    FSM_sub_bytes_0_t110 = 64'b0000000000000000000000000000000000000000000000000000000000001010;
    FSM_sub_bytes_0_t111 = FSM_sub_bytes_0_t110[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t112 = 64'b0000000000000000000000000000000000000000000000000000000000001010;
    FSM_sub_bytes_0_t113 = FSM_sub_bytes_0_t112[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t114 = FSM_sub_bytes_0_t109[FSM_sub_bytes_0_t113 * 64 +: 64];
    FSM_sub_bytes_0_t115 = FSM_sub_bytes_0_t114[6'b0 * 1 +: 8 * 1];
    FSM_sub_bytes_0_t116 = FSM_sub_bytes_0_t31[FSM_sub_bytes_0_t115 * 64 +: 64];
    FSM_sub_bytes_0_t117 = FSM_sub_bytes_0_t109;
    FSM_sub_bytes_0_t117[FSM_sub_bytes_0_t111 * 64 +: 64] = FSM_sub_bytes_0_t116;
    FSM_sub_bytes_0_t118 = 64'b0000000000000000000000000000000000000000000000000000000000001011;
    FSM_sub_bytes_0_t119 = FSM_sub_bytes_0_t118[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t120 = 64'b0000000000000000000000000000000000000000000000000000000000001011;
    FSM_sub_bytes_0_t121 = FSM_sub_bytes_0_t120[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t122 = FSM_sub_bytes_0_t117[FSM_sub_bytes_0_t121 * 64 +: 64];
    FSM_sub_bytes_0_t123 = FSM_sub_bytes_0_t122[6'b0 * 1 +: 8 * 1];
    FSM_sub_bytes_0_t124 = FSM_sub_bytes_0_t31[FSM_sub_bytes_0_t123 * 64 +: 64];
    FSM_sub_bytes_0_t125 = FSM_sub_bytes_0_t117;
    FSM_sub_bytes_0_t125[FSM_sub_bytes_0_t119 * 64 +: 64] = FSM_sub_bytes_0_t124;
    FSM_sub_bytes_0_t126 = 64'b0000000000000000000000000000000000000000000000000000000000001100;
    FSM_sub_bytes_0_t127 = FSM_sub_bytes_0_t126[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t128 = 64'b0000000000000000000000000000000000000000000000000000000000001100;
    FSM_sub_bytes_0_t129 = FSM_sub_bytes_0_t128[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t130 = FSM_sub_bytes_0_t125[FSM_sub_bytes_0_t129 * 64 +: 64];
    FSM_sub_bytes_0_t131 = FSM_sub_bytes_0_t130[6'b0 * 1 +: 8 * 1];
    FSM_sub_bytes_0_t132 = FSM_sub_bytes_0_t31[FSM_sub_bytes_0_t131 * 64 +: 64];
    FSM_sub_bytes_0_t133 = FSM_sub_bytes_0_t125;
    FSM_sub_bytes_0_t133[FSM_sub_bytes_0_t127 * 64 +: 64] = FSM_sub_bytes_0_t132;
    FSM_sub_bytes_0_t134 = 64'b0000000000000000000000000000000000000000000000000000000000001101;
    FSM_sub_bytes_0_t135 = FSM_sub_bytes_0_t134[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t136 = 64'b0000000000000000000000000000000000000000000000000000000000001101;
    FSM_sub_bytes_0_t137 = FSM_sub_bytes_0_t136[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t138 = FSM_sub_bytes_0_t133[FSM_sub_bytes_0_t137 * 64 +: 64];
    FSM_sub_bytes_0_t139 = FSM_sub_bytes_0_t138[6'b0 * 1 +: 8 * 1];
    FSM_sub_bytes_0_t140 = FSM_sub_bytes_0_t31[FSM_sub_bytes_0_t139 * 64 +: 64];
    FSM_sub_bytes_0_t141 = FSM_sub_bytes_0_t133;
    FSM_sub_bytes_0_t141[FSM_sub_bytes_0_t135 * 64 +: 64] = FSM_sub_bytes_0_t140;
    FSM_sub_bytes_0_t142 = 64'b0000000000000000000000000000000000000000000000000000000000001110;
    FSM_sub_bytes_0_t143 = FSM_sub_bytes_0_t142[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t144 = 64'b0000000000000000000000000000000000000000000000000000000000001110;
    FSM_sub_bytes_0_t145 = FSM_sub_bytes_0_t144[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t146 = FSM_sub_bytes_0_t141[FSM_sub_bytes_0_t145 * 64 +: 64];
    FSM_sub_bytes_0_t147 = FSM_sub_bytes_0_t146[6'b0 * 1 +: 8 * 1];
    FSM_sub_bytes_0_t148 = FSM_sub_bytes_0_t31[FSM_sub_bytes_0_t147 * 64 +: 64];
    FSM_sub_bytes_0_t149 = FSM_sub_bytes_0_t141;
    FSM_sub_bytes_0_t149[FSM_sub_bytes_0_t143 * 64 +: 64] = FSM_sub_bytes_0_t148;
    FSM_sub_bytes_0_t150 = 64'b0000000000000000000000000000000000000000000000000000000000001111;
    FSM_sub_bytes_0_t151 = FSM_sub_bytes_0_t150[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t152 = 64'b0000000000000000000000000000000000000000000000000000000000001111;
    FSM_sub_bytes_0_t153 = FSM_sub_bytes_0_t152[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t154 = FSM_sub_bytes_0_t149[FSM_sub_bytes_0_t153 * 64 +: 64];
    FSM_sub_bytes_0_t155 = FSM_sub_bytes_0_t154[6'b0 * 1 +: 8 * 1];
    FSM_sub_bytes_0_t156 = FSM_sub_bytes_0_t31[FSM_sub_bytes_0_t155 * 64 +: 64];
    FSM_sub_bytes_0_t157 = FSM_sub_bytes_0_t149;
    FSM_sub_bytes_0_t157[FSM_sub_bytes_0_t151 * 64 +: 64] = FSM_sub_bytes_0_t156;
    FSM_sub_bytes_0_t158 = 64'b0;
    FSM_sub_bytes_0_t159 = FSM_sub_bytes_0_t158[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t160 = FSM_sub_bytes_0_t157[FSM_sub_bytes_0_t159 * 64 +: 64];
    FSM_sub_bytes_0_t161 = 64'b0000000000000000000000000000000000000000000000000000000000000001;
    FSM_sub_bytes_0_t162 = FSM_sub_bytes_0_t161[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t163 = FSM_sub_bytes_0_t157[FSM_sub_bytes_0_t162 * 64 +: 64];
    FSM_sub_bytes_0_t164 = 64'b0000000000000000000000000000000000000000000000000000000000001000;
    FSM_sub_bytes_0_t165 = FSM_sub_bytes_0_t164[6'b0 * 1 +: 6 * 1];
    FSM_sub_bytes_0_t166 = 64'b0000000000000000000000000000000000000000000000000000000000000010;
    FSM_sub_bytes_0_t167 = FSM_sub_bytes_0_t166[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t168 = FSM_sub_bytes_0_t157[FSM_sub_bytes_0_t167 * 64 +: 64];
    FSM_sub_bytes_0_t169 = 64'b0000000000000000000000000000000000000000000000000000000000010000;
    FSM_sub_bytes_0_t170 = FSM_sub_bytes_0_t169[6'b0 * 1 +: 6 * 1];
    FSM_sub_bytes_0_t171 = 64'b0000000000000000000000000000000000000000000000000000000000000011;
    FSM_sub_bytes_0_t172 = FSM_sub_bytes_0_t171[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t173 = FSM_sub_bytes_0_t157[FSM_sub_bytes_0_t172 * 64 +: 64];
    FSM_sub_bytes_0_t174 = 64'b0000000000000000000000000000000000000000000000000000000000011000;
    FSM_sub_bytes_0_t175 = FSM_sub_bytes_0_t174[6'b0 * 1 +: 6 * 1];
    FSM_sub_bytes_0_t176 = 64'b0000000000000000000000000000000000000000000000000000000000000100;
    FSM_sub_bytes_0_t177 = FSM_sub_bytes_0_t176[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t178 = FSM_sub_bytes_0_t157[FSM_sub_bytes_0_t177 * 64 +: 64];
    FSM_sub_bytes_0_t179 = 64'b0000000000000000000000000000000000000000000000000000000000100000;
    FSM_sub_bytes_0_t180 = FSM_sub_bytes_0_t179[6'b0 * 1 +: 6 * 1];
    FSM_sub_bytes_0_t181 = 64'b0000000000000000000000000000000000000000000000000000000000000101;
    FSM_sub_bytes_0_t182 = FSM_sub_bytes_0_t181[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t183 = FSM_sub_bytes_0_t157[FSM_sub_bytes_0_t182 * 64 +: 64];
    FSM_sub_bytes_0_t184 = 64'b0000000000000000000000000000000000000000000000000000000000101000;
    FSM_sub_bytes_0_t185 = FSM_sub_bytes_0_t184[6'b0 * 1 +: 6 * 1];
    FSM_sub_bytes_0_t186 = 64'b0000000000000000000000000000000000000000000000000000000000000110;
    FSM_sub_bytes_0_t187 = FSM_sub_bytes_0_t186[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t188 = FSM_sub_bytes_0_t157[FSM_sub_bytes_0_t187 * 64 +: 64];
    FSM_sub_bytes_0_t189 = 64'b0000000000000000000000000000000000000000000000000000000000110000;
    FSM_sub_bytes_0_t190 = FSM_sub_bytes_0_t189[6'b0 * 1 +: 6 * 1];
    FSM_sub_bytes_0_t191 = 64'b0000000000000000000000000000000000000000000000000000000000000111;
    FSM_sub_bytes_0_t192 = FSM_sub_bytes_0_t191[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t193 = FSM_sub_bytes_0_t157[FSM_sub_bytes_0_t192 * 64 +: 64];
    FSM_sub_bytes_0_t194 = 64'b0000000000000000000000000000000000000000000000000000000000111000;
    FSM_sub_bytes_0_t195 = FSM_sub_bytes_0_t194[6'b0 * 1 +: 6 * 1];
    FSM_sub_bytes_0_t196 = 64'b0000000000000000000000000000000000000000000000000000000000001000;
    FSM_sub_bytes_0_t197 = FSM_sub_bytes_0_t196[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t198 = FSM_sub_bytes_0_t157[FSM_sub_bytes_0_t197 * 64 +: 64];
    FSM_sub_bytes_0_t199 = 64'b0000000000000000000000000000000000000000000000000000000000001001;
    FSM_sub_bytes_0_t200 = FSM_sub_bytes_0_t199[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t201 = FSM_sub_bytes_0_t157[FSM_sub_bytes_0_t200 * 64 +: 64];
    FSM_sub_bytes_0_t202 = 64'b0000000000000000000000000000000000000000000000000000000000001000;
    FSM_sub_bytes_0_t203 = FSM_sub_bytes_0_t202[6'b0 * 1 +: 6 * 1];
    FSM_sub_bytes_0_t204 = 64'b0000000000000000000000000000000000000000000000000000000000001010;
    FSM_sub_bytes_0_t205 = FSM_sub_bytes_0_t204[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t206 = FSM_sub_bytes_0_t157[FSM_sub_bytes_0_t205 * 64 +: 64];
    FSM_sub_bytes_0_t207 = 64'b0000000000000000000000000000000000000000000000000000000000010000;
    FSM_sub_bytes_0_t208 = FSM_sub_bytes_0_t207[6'b0 * 1 +: 6 * 1];
    FSM_sub_bytes_0_t209 = 64'b0000000000000000000000000000000000000000000000000000000000001011;
    FSM_sub_bytes_0_t210 = FSM_sub_bytes_0_t209[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t211 = FSM_sub_bytes_0_t157[FSM_sub_bytes_0_t210 * 64 +: 64];
    FSM_sub_bytes_0_t212 = 64'b0000000000000000000000000000000000000000000000000000000000011000;
    FSM_sub_bytes_0_t213 = FSM_sub_bytes_0_t212[6'b0 * 1 +: 6 * 1];
    FSM_sub_bytes_0_t214 = 64'b0000000000000000000000000000000000000000000000000000000000001100;
    FSM_sub_bytes_0_t215 = FSM_sub_bytes_0_t214[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t216 = FSM_sub_bytes_0_t157[FSM_sub_bytes_0_t215 * 64 +: 64];
    FSM_sub_bytes_0_t217 = 64'b0000000000000000000000000000000000000000000000000000000000100000;
    FSM_sub_bytes_0_t218 = FSM_sub_bytes_0_t217[6'b0 * 1 +: 6 * 1];
    FSM_sub_bytes_0_t219 = 64'b0000000000000000000000000000000000000000000000000000000000001101;
    FSM_sub_bytes_0_t220 = FSM_sub_bytes_0_t219[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t221 = FSM_sub_bytes_0_t157[FSM_sub_bytes_0_t220 * 64 +: 64];
    FSM_sub_bytes_0_t222 = 64'b0000000000000000000000000000000000000000000000000000000000101000;
    FSM_sub_bytes_0_t223 = FSM_sub_bytes_0_t222[6'b0 * 1 +: 6 * 1];
    FSM_sub_bytes_0_t224 = 64'b0000000000000000000000000000000000000000000000000000000000001110;
    FSM_sub_bytes_0_t225 = FSM_sub_bytes_0_t224[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t226 = FSM_sub_bytes_0_t157[FSM_sub_bytes_0_t225 * 64 +: 64];
    FSM_sub_bytes_0_t227 = 64'b0000000000000000000000000000000000000000000000000000000000110000;
    FSM_sub_bytes_0_t228 = FSM_sub_bytes_0_t227[6'b0 * 1 +: 6 * 1];
    FSM_sub_bytes_0_t229 = 64'b0000000000000000000000000000000000000000000000000000000000001111;
    FSM_sub_bytes_0_t230 = FSM_sub_bytes_0_t229[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t231 = FSM_sub_bytes_0_t157[FSM_sub_bytes_0_t230 * 64 +: 64];
    FSM_sub_bytes_0_t232 = 64'b0000000000000000000000000000000000000000000000000000000000111000;
    FSM_sub_bytes_0_t233 = FSM_sub_bytes_0_t232[6'b0 * 1 +: 6 * 1];
end

always @* begin
    FSM_sub_bytes_0_t0[0 * 64 +: 64] = i_lower_bits & 64'b0000000000000000000000000000000000000000000000000000000011111111;
    FSM_sub_bytes_0_t1 = 64'b0000000000000000000000000000000000000000000000000000000000001000;
    FSM_sub_bytes_0_t2 = FSM_sub_bytes_0_t1[6'b0 * 1 +: 6 * 1];
    FSM_sub_bytes_0_t0[1 * 64 +: 64] = (i_lower_bits >> FSM_sub_bytes_0_t2) & 64'b0000000000000000000000000000000000000000000000000000000011111111;
    FSM_sub_bytes_0_t3 = 64'b0000000000000000000000000000000000000000000000000000000000010000;
    FSM_sub_bytes_0_t4 = FSM_sub_bytes_0_t3[6'b0 * 1 +: 6 * 1];
    FSM_sub_bytes_0_t0[2 * 64 +: 64] = (i_lower_bits >> FSM_sub_bytes_0_t4) & 64'b0000000000000000000000000000000000000000000000000000000011111111;
    FSM_sub_bytes_0_t5 = 64'b0000000000000000000000000000000000000000000000000000000000011000;
    FSM_sub_bytes_0_t6 = FSM_sub_bytes_0_t5[6'b0 * 1 +: 6 * 1];
    FSM_sub_bytes_0_t0[3 * 64 +: 64] = (i_lower_bits >> FSM_sub_bytes_0_t6) & 64'b0000000000000000000000000000000000000000000000000000000011111111;
    FSM_sub_bytes_0_t7 = 64'b0000000000000000000000000000000000000000000000000000000000100000;
    FSM_sub_bytes_0_t8 = FSM_sub_bytes_0_t7[6'b0 * 1 +: 6 * 1];
    FSM_sub_bytes_0_t0[4 * 64 +: 64] = (i_lower_bits >> FSM_sub_bytes_0_t8) & 64'b0000000000000000000000000000000000000000000000000000000011111111;
    FSM_sub_bytes_0_t9 = 64'b0000000000000000000000000000000000000000000000000000000000101000;
    FSM_sub_bytes_0_t10 = FSM_sub_bytes_0_t9[6'b0 * 1 +: 6 * 1];
    FSM_sub_bytes_0_t0[5 * 64 +: 64] = (i_lower_bits >> FSM_sub_bytes_0_t10) & 64'b0000000000000000000000000000000000000000000000000000000011111111;
    FSM_sub_bytes_0_t11 = 64'b0000000000000000000000000000000000000000000000000000000000110000;
    FSM_sub_bytes_0_t12 = FSM_sub_bytes_0_t11[6'b0 * 1 +: 6 * 1];
    FSM_sub_bytes_0_t0[6 * 64 +: 64] = (i_lower_bits >> FSM_sub_bytes_0_t12) & 64'b0000000000000000000000000000000000000000000000000000000011111111;
    FSM_sub_bytes_0_t13 = 64'b0000000000000000000000000000000000000000000000000000000000111000;
    FSM_sub_bytes_0_t14 = FSM_sub_bytes_0_t13[6'b0 * 1 +: 6 * 1];
    FSM_sub_bytes_0_t0[7 * 64 +: 64] = (i_lower_bits >> FSM_sub_bytes_0_t14) & 64'b0000000000000000000000000000000000000000000000000000000011111111;
    FSM_sub_bytes_0_t0[8 * 64 +: 64] = i_higher_bits & 64'b0000000000000000000000000000000000000000000000000000000011111111;
    FSM_sub_bytes_0_t15 = 64'b0000000000000000000000000000000000000000000000000000000000001000;
    FSM_sub_bytes_0_t16 = FSM_sub_bytes_0_t15[6'b0 * 1 +: 6 * 1];
    FSM_sub_bytes_0_t0[9 * 64 +: 64] = (i_higher_bits >> FSM_sub_bytes_0_t16) & 64'b0000000000000000000000000000000000000000000000000000000011111111;
    FSM_sub_bytes_0_t17 = 64'b0000000000000000000000000000000000000000000000000000000000010000;
    FSM_sub_bytes_0_t18 = FSM_sub_bytes_0_t17[6'b0 * 1 +: 6 * 1];
    FSM_sub_bytes_0_t0[10 * 64 +: 64] = (i_higher_bits >> FSM_sub_bytes_0_t18) & 64'b0000000000000000000000000000000000000000000000000000000011111111;
    FSM_sub_bytes_0_t19 = 64'b0000000000000000000000000000000000000000000000000000000000011000;
    FSM_sub_bytes_0_t20 = FSM_sub_bytes_0_t19[6'b0 * 1 +: 6 * 1];
    FSM_sub_bytes_0_t0[11 * 64 +: 64] = (i_higher_bits >> FSM_sub_bytes_0_t20) & 64'b0000000000000000000000000000000000000000000000000000000011111111;
    FSM_sub_bytes_0_t21 = 64'b0000000000000000000000000000000000000000000000000000000000100000;
    FSM_sub_bytes_0_t22 = FSM_sub_bytes_0_t21[6'b0 * 1 +: 6 * 1];
    FSM_sub_bytes_0_t0[12 * 64 +: 64] = (i_higher_bits >> FSM_sub_bytes_0_t22) & 64'b0000000000000000000000000000000000000000000000000000000011111111;
    FSM_sub_bytes_0_t23 = 64'b0000000000000000000000000000000000000000000000000000000000101000;
    FSM_sub_bytes_0_t24 = FSM_sub_bytes_0_t23[6'b0 * 1 +: 6 * 1];
    FSM_sub_bytes_0_t0[13 * 64 +: 64] = (i_higher_bits >> FSM_sub_bytes_0_t24) & 64'b0000000000000000000000000000000000000000000000000000000011111111;
    FSM_sub_bytes_0_t25 = 64'b0000000000000000000000000000000000000000000000000000000000110000;
    FSM_sub_bytes_0_t26 = FSM_sub_bytes_0_t25[6'b0 * 1 +: 6 * 1];
    FSM_sub_bytes_0_t0[14 * 64 +: 64] = (i_higher_bits >> FSM_sub_bytes_0_t26) & 64'b0000000000000000000000000000000000000000000000000000000011111111;
    FSM_sub_bytes_0_t27 = 64'b0000000000000000000000000000000000000000000000000000000000111000;
    FSM_sub_bytes_0_t28 = FSM_sub_bytes_0_t27[6'b0 * 1 +: 6 * 1];
    FSM_sub_bytes_0_t0[15 * 64 +: 64] = (i_higher_bits >> FSM_sub_bytes_0_t28) & 64'b0000000000000000000000000000000000000000000000000000000011111111;
    FSM_sub_bytes_0_t29 = 64'b0;
    FSM_sub_bytes_0_t30 = FSM_sub_bytes_0_t29[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t31[0 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001100011;
    FSM_sub_bytes_0_t31[1 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001111100;
    FSM_sub_bytes_0_t31[2 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001110111;
    FSM_sub_bytes_0_t31[3 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001111011;
    FSM_sub_bytes_0_t31[4 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011110010;
    FSM_sub_bytes_0_t31[5 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001101011;
    FSM_sub_bytes_0_t31[6 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001101111;
    FSM_sub_bytes_0_t31[7 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011000101;
    FSM_sub_bytes_0_t31[8 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000110000;
    FSM_sub_bytes_0_t31[9 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000000001;
    FSM_sub_bytes_0_t31[10 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001100111;
    FSM_sub_bytes_0_t31[11 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000101011;
    FSM_sub_bytes_0_t31[12 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011111110;
    FSM_sub_bytes_0_t31[13 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011010111;
    FSM_sub_bytes_0_t31[14 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010101011;
    FSM_sub_bytes_0_t31[15 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001110110;
    FSM_sub_bytes_0_t31[16 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011001010;
    FSM_sub_bytes_0_t31[17 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010000010;
    FSM_sub_bytes_0_t31[18 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011001001;
    FSM_sub_bytes_0_t31[19 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001111101;
    FSM_sub_bytes_0_t31[20 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011111010;
    FSM_sub_bytes_0_t31[21 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001011001;
    FSM_sub_bytes_0_t31[22 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001000111;
    FSM_sub_bytes_0_t31[23 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011110000;
    FSM_sub_bytes_0_t31[24 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010101101;
    FSM_sub_bytes_0_t31[25 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011010100;
    FSM_sub_bytes_0_t31[26 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010100010;
    FSM_sub_bytes_0_t31[27 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010101111;
    FSM_sub_bytes_0_t31[28 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010011100;
    FSM_sub_bytes_0_t31[29 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010100100;
    FSM_sub_bytes_0_t31[30 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001110010;
    FSM_sub_bytes_0_t31[31 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011000000;
    FSM_sub_bytes_0_t31[32 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010110111;
    FSM_sub_bytes_0_t31[33 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011111101;
    FSM_sub_bytes_0_t31[34 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010010011;
    FSM_sub_bytes_0_t31[35 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000100110;
    FSM_sub_bytes_0_t31[36 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000110110;
    FSM_sub_bytes_0_t31[37 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000111111;
    FSM_sub_bytes_0_t31[38 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011110111;
    FSM_sub_bytes_0_t31[39 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011001100;
    FSM_sub_bytes_0_t31[40 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000110100;
    FSM_sub_bytes_0_t31[41 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010100101;
    FSM_sub_bytes_0_t31[42 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011100101;
    FSM_sub_bytes_0_t31[43 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011110001;
    FSM_sub_bytes_0_t31[44 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001110001;
    FSM_sub_bytes_0_t31[45 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011011000;
    FSM_sub_bytes_0_t31[46 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000110001;
    FSM_sub_bytes_0_t31[47 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000010101;
    FSM_sub_bytes_0_t31[48 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000000100;
    FSM_sub_bytes_0_t31[49 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011000111;
    FSM_sub_bytes_0_t31[50 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000100011;
    FSM_sub_bytes_0_t31[51 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011000011;
    FSM_sub_bytes_0_t31[52 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000011000;
    FSM_sub_bytes_0_t31[53 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010010110;
    FSM_sub_bytes_0_t31[54 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000000101;
    FSM_sub_bytes_0_t31[55 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010011010;
    FSM_sub_bytes_0_t31[56 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000000111;
    FSM_sub_bytes_0_t31[57 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000010010;
    FSM_sub_bytes_0_t31[58 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010000000;
    FSM_sub_bytes_0_t31[59 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011100010;
    FSM_sub_bytes_0_t31[60 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011101011;
    FSM_sub_bytes_0_t31[61 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000100111;
    FSM_sub_bytes_0_t31[62 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010110010;
    FSM_sub_bytes_0_t31[63 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001110101;
    FSM_sub_bytes_0_t31[64 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000001001;
    FSM_sub_bytes_0_t31[65 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010000011;
    FSM_sub_bytes_0_t31[66 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000101100;
    FSM_sub_bytes_0_t31[67 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000011010;
    FSM_sub_bytes_0_t31[68 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000011011;
    FSM_sub_bytes_0_t31[69 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001101110;
    FSM_sub_bytes_0_t31[70 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001011010;
    FSM_sub_bytes_0_t31[71 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010100000;
    FSM_sub_bytes_0_t31[72 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001010010;
    FSM_sub_bytes_0_t31[73 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000111011;
    FSM_sub_bytes_0_t31[74 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011010110;
    FSM_sub_bytes_0_t31[75 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010110011;
    FSM_sub_bytes_0_t31[76 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000101001;
    FSM_sub_bytes_0_t31[77 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011100011;
    FSM_sub_bytes_0_t31[78 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000101111;
    FSM_sub_bytes_0_t31[79 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010000100;
    FSM_sub_bytes_0_t31[80 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001010011;
    FSM_sub_bytes_0_t31[81 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011010001;
    FSM_sub_bytes_0_t31[82 * 64 +: 64] = 64'b0;
    FSM_sub_bytes_0_t31[83 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011101101;
    FSM_sub_bytes_0_t31[84 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000100000;
    FSM_sub_bytes_0_t31[85 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011111100;
    FSM_sub_bytes_0_t31[86 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010110001;
    FSM_sub_bytes_0_t31[87 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001011011;
    FSM_sub_bytes_0_t31[88 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001101010;
    FSM_sub_bytes_0_t31[89 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011001011;
    FSM_sub_bytes_0_t31[90 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010111110;
    FSM_sub_bytes_0_t31[91 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000111001;
    FSM_sub_bytes_0_t31[92 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001001010;
    FSM_sub_bytes_0_t31[93 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001001100;
    FSM_sub_bytes_0_t31[94 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001011000;
    FSM_sub_bytes_0_t31[95 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011001111;
    FSM_sub_bytes_0_t31[96 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011010000;
    FSM_sub_bytes_0_t31[97 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011101111;
    FSM_sub_bytes_0_t31[98 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010101010;
    FSM_sub_bytes_0_t31[99 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011111011;
    FSM_sub_bytes_0_t31[100 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001000011;
    FSM_sub_bytes_0_t31[101 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001001101;
    FSM_sub_bytes_0_t31[102 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000110011;
    FSM_sub_bytes_0_t31[103 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010000101;
    FSM_sub_bytes_0_t31[104 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001000101;
    FSM_sub_bytes_0_t31[105 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011111001;
    FSM_sub_bytes_0_t31[106 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000000010;
    FSM_sub_bytes_0_t31[107 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001111111;
    FSM_sub_bytes_0_t31[108 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001010000;
    FSM_sub_bytes_0_t31[109 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000111100;
    FSM_sub_bytes_0_t31[110 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010011111;
    FSM_sub_bytes_0_t31[111 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010101000;
    FSM_sub_bytes_0_t31[112 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001010001;
    FSM_sub_bytes_0_t31[113 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010100011;
    FSM_sub_bytes_0_t31[114 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001000000;
    FSM_sub_bytes_0_t31[115 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010001111;
    FSM_sub_bytes_0_t31[116 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010010010;
    FSM_sub_bytes_0_t31[117 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010011101;
    FSM_sub_bytes_0_t31[118 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000111000;
    FSM_sub_bytes_0_t31[119 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011110101;
    FSM_sub_bytes_0_t31[120 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010111100;
    FSM_sub_bytes_0_t31[121 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010110110;
    FSM_sub_bytes_0_t31[122 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011011010;
    FSM_sub_bytes_0_t31[123 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000100001;
    FSM_sub_bytes_0_t31[124 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000010000;
    FSM_sub_bytes_0_t31[125 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011111111;
    FSM_sub_bytes_0_t31[126 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011110011;
    FSM_sub_bytes_0_t31[127 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011010010;
    FSM_sub_bytes_0_t31[128 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011001101;
    FSM_sub_bytes_0_t31[129 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000001100;
    FSM_sub_bytes_0_t31[130 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000010011;
    FSM_sub_bytes_0_t31[131 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011101100;
    FSM_sub_bytes_0_t31[132 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001011111;
    FSM_sub_bytes_0_t31[133 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010010111;
    FSM_sub_bytes_0_t31[134 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001000100;
    FSM_sub_bytes_0_t31[135 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000010111;
    FSM_sub_bytes_0_t31[136 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011000100;
    FSM_sub_bytes_0_t31[137 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010100111;
    FSM_sub_bytes_0_t31[138 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001111110;
    FSM_sub_bytes_0_t31[139 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000111101;
    FSM_sub_bytes_0_t31[140 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001100100;
    FSM_sub_bytes_0_t31[141 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001011101;
    FSM_sub_bytes_0_t31[142 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000011001;
    FSM_sub_bytes_0_t31[143 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001110011;
    FSM_sub_bytes_0_t31[144 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001100000;
    FSM_sub_bytes_0_t31[145 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010000001;
    FSM_sub_bytes_0_t31[146 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001001111;
    FSM_sub_bytes_0_t31[147 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011011100;
    FSM_sub_bytes_0_t31[148 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000100010;
    FSM_sub_bytes_0_t31[149 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000101010;
    FSM_sub_bytes_0_t31[150 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010010000;
    FSM_sub_bytes_0_t31[151 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010001000;
    FSM_sub_bytes_0_t31[152 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001000110;
    FSM_sub_bytes_0_t31[153 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011101110;
    FSM_sub_bytes_0_t31[154 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010111000;
    FSM_sub_bytes_0_t31[155 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000010100;
    FSM_sub_bytes_0_t31[156 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011011110;
    FSM_sub_bytes_0_t31[157 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001011110;
    FSM_sub_bytes_0_t31[158 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000001011;
    FSM_sub_bytes_0_t31[159 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011011011;
    FSM_sub_bytes_0_t31[160 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011100000;
    FSM_sub_bytes_0_t31[161 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000110010;
    FSM_sub_bytes_0_t31[162 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000111010;
    FSM_sub_bytes_0_t31[163 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000001010;
    FSM_sub_bytes_0_t31[164 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001001001;
    FSM_sub_bytes_0_t31[165 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000000110;
    FSM_sub_bytes_0_t31[166 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000100100;
    FSM_sub_bytes_0_t31[167 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001011100;
    FSM_sub_bytes_0_t31[168 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011000010;
    FSM_sub_bytes_0_t31[169 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011010011;
    FSM_sub_bytes_0_t31[170 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010101100;
    FSM_sub_bytes_0_t31[171 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001100010;
    FSM_sub_bytes_0_t31[172 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010010001;
    FSM_sub_bytes_0_t31[173 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010010101;
    FSM_sub_bytes_0_t31[174 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011100100;
    FSM_sub_bytes_0_t31[175 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001111001;
    FSM_sub_bytes_0_t31[176 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011100111;
    FSM_sub_bytes_0_t31[177 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011001000;
    FSM_sub_bytes_0_t31[178 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000110111;
    FSM_sub_bytes_0_t31[179 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001101101;
    FSM_sub_bytes_0_t31[180 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010001101;
    FSM_sub_bytes_0_t31[181 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011010101;
    FSM_sub_bytes_0_t31[182 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001001110;
    FSM_sub_bytes_0_t31[183 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010101001;
    FSM_sub_bytes_0_t31[184 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001101100;
    FSM_sub_bytes_0_t31[185 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001010110;
    FSM_sub_bytes_0_t31[186 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011110100;
    FSM_sub_bytes_0_t31[187 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011101010;
    FSM_sub_bytes_0_t31[188 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001100101;
    FSM_sub_bytes_0_t31[189 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001111010;
    FSM_sub_bytes_0_t31[190 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010101110;
    FSM_sub_bytes_0_t31[191 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000001000;
    FSM_sub_bytes_0_t31[192 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010111010;
    FSM_sub_bytes_0_t31[193 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001111000;
    FSM_sub_bytes_0_t31[194 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000100101;
    FSM_sub_bytes_0_t31[195 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000101110;
    FSM_sub_bytes_0_t31[196 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000011100;
    FSM_sub_bytes_0_t31[197 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010100110;
    FSM_sub_bytes_0_t31[198 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010110100;
    FSM_sub_bytes_0_t31[199 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011000110;
    FSM_sub_bytes_0_t31[200 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011101000;
    FSM_sub_bytes_0_t31[201 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011011101;
    FSM_sub_bytes_0_t31[202 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001110100;
    FSM_sub_bytes_0_t31[203 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000011111;
    FSM_sub_bytes_0_t31[204 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001001011;
    FSM_sub_bytes_0_t31[205 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010111101;
    FSM_sub_bytes_0_t31[206 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010001011;
    FSM_sub_bytes_0_t31[207 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010001010;
    FSM_sub_bytes_0_t31[208 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001110000;
    FSM_sub_bytes_0_t31[209 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000111110;
    FSM_sub_bytes_0_t31[210 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010110101;
    FSM_sub_bytes_0_t31[211 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001100110;
    FSM_sub_bytes_0_t31[212 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001001000;
    FSM_sub_bytes_0_t31[213 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000000011;
    FSM_sub_bytes_0_t31[214 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011110110;
    FSM_sub_bytes_0_t31[215 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000001110;
    FSM_sub_bytes_0_t31[216 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001100001;
    FSM_sub_bytes_0_t31[217 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000110101;
    FSM_sub_bytes_0_t31[218 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001010111;
    FSM_sub_bytes_0_t31[219 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010111001;
    FSM_sub_bytes_0_t31[220 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010000110;
    FSM_sub_bytes_0_t31[221 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011000001;
    FSM_sub_bytes_0_t31[222 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000011101;
    FSM_sub_bytes_0_t31[223 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010011110;
    FSM_sub_bytes_0_t31[224 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011100001;
    FSM_sub_bytes_0_t31[225 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011111000;
    FSM_sub_bytes_0_t31[226 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010011000;
    FSM_sub_bytes_0_t31[227 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000010001;
    FSM_sub_bytes_0_t31[228 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001101001;
    FSM_sub_bytes_0_t31[229 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011011001;
    FSM_sub_bytes_0_t31[230 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010001110;
    FSM_sub_bytes_0_t31[231 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010010100;
    FSM_sub_bytes_0_t31[232 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010011011;
    FSM_sub_bytes_0_t31[233 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000011110;
    FSM_sub_bytes_0_t31[234 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010000111;
    FSM_sub_bytes_0_t31[235 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011101001;
    FSM_sub_bytes_0_t31[236 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011001110;
    FSM_sub_bytes_0_t31[237 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001010101;
    FSM_sub_bytes_0_t31[238 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000101000;
    FSM_sub_bytes_0_t31[239 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011011111;
    FSM_sub_bytes_0_t31[240 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010001100;
    FSM_sub_bytes_0_t31[241 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010100001;
    FSM_sub_bytes_0_t31[242 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010001001;
    FSM_sub_bytes_0_t31[243 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000001101;
    FSM_sub_bytes_0_t31[244 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010111111;
    FSM_sub_bytes_0_t31[245 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000011100110;
    FSM_sub_bytes_0_t31[246 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001000010;
    FSM_sub_bytes_0_t31[247 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001101000;
    FSM_sub_bytes_0_t31[248 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001000001;
    FSM_sub_bytes_0_t31[249 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010011001;
    FSM_sub_bytes_0_t31[250 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000101101;
    FSM_sub_bytes_0_t31[251 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000001111;
    FSM_sub_bytes_0_t31[252 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010110000;
    FSM_sub_bytes_0_t31[253 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000001010100;
    FSM_sub_bytes_0_t31[254 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000010111011;
    FSM_sub_bytes_0_t31[255 * 64 +: 64] = 64'b0000000000000000000000000000000000000000000000000000000000010110;
    FSM_sub_bytes_0_t32 = 64'b0;
    FSM_sub_bytes_0_t33 = FSM_sub_bytes_0_t32[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t34 = FSM_sub_bytes_0_t0[FSM_sub_bytes_0_t33 * 64 +: 64];
    FSM_sub_bytes_0_t35 = FSM_sub_bytes_0_t34[6'b0 * 1 +: 8 * 1];
    FSM_sub_bytes_0_t36 = FSM_sub_bytes_0_t31[FSM_sub_bytes_0_t35 * 64 +: 64];
    FSM_sub_bytes_0_t37 = FSM_sub_bytes_0_t0;
    FSM_sub_bytes_0_t37[FSM_sub_bytes_0_t30 * 64 +: 64] = FSM_sub_bytes_0_t36;
    FSM_sub_bytes_0_t38 = 64'b0000000000000000000000000000000000000000000000000000000000000001;
    FSM_sub_bytes_0_t39 = FSM_sub_bytes_0_t38[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t40 = 64'b0000000000000000000000000000000000000000000000000000000000000001;
    FSM_sub_bytes_0_t41 = FSM_sub_bytes_0_t40[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t42 = FSM_sub_bytes_0_t37[FSM_sub_bytes_0_t41 * 64 +: 64];
    FSM_sub_bytes_0_t43 = FSM_sub_bytes_0_t42[6'b0 * 1 +: 8 * 1];
    FSM_sub_bytes_0_t44 = FSM_sub_bytes_0_t31[FSM_sub_bytes_0_t43 * 64 +: 64];
    FSM_sub_bytes_0_t45 = FSM_sub_bytes_0_t37;
    FSM_sub_bytes_0_t45[FSM_sub_bytes_0_t39 * 64 +: 64] = FSM_sub_bytes_0_t44;
    FSM_sub_bytes_0_t46 = 64'b0000000000000000000000000000000000000000000000000000000000000010;
    FSM_sub_bytes_0_t47 = FSM_sub_bytes_0_t46[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t48 = 64'b0000000000000000000000000000000000000000000000000000000000000010;
    FSM_sub_bytes_0_t49 = FSM_sub_bytes_0_t48[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t50 = FSM_sub_bytes_0_t45[FSM_sub_bytes_0_t49 * 64 +: 64];
    FSM_sub_bytes_0_t51 = FSM_sub_bytes_0_t50[6'b0 * 1 +: 8 * 1];
    FSM_sub_bytes_0_t52 = FSM_sub_bytes_0_t31[FSM_sub_bytes_0_t51 * 64 +: 64];
    FSM_sub_bytes_0_t53 = FSM_sub_bytes_0_t45;
    FSM_sub_bytes_0_t53[FSM_sub_bytes_0_t47 * 64 +: 64] = FSM_sub_bytes_0_t52;
    FSM_sub_bytes_0_t54 = 64'b0000000000000000000000000000000000000000000000000000000000000011;
    FSM_sub_bytes_0_t55 = FSM_sub_bytes_0_t54[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t56 = 64'b0000000000000000000000000000000000000000000000000000000000000011;
    FSM_sub_bytes_0_t57 = FSM_sub_bytes_0_t56[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t58 = FSM_sub_bytes_0_t53[FSM_sub_bytes_0_t57 * 64 +: 64];
    FSM_sub_bytes_0_t59 = FSM_sub_bytes_0_t58[6'b0 * 1 +: 8 * 1];
    FSM_sub_bytes_0_t60 = FSM_sub_bytes_0_t31[FSM_sub_bytes_0_t59 * 64 +: 64];
    FSM_sub_bytes_0_t61 = FSM_sub_bytes_0_t53;
    FSM_sub_bytes_0_t61[FSM_sub_bytes_0_t55 * 64 +: 64] = FSM_sub_bytes_0_t60;
    FSM_sub_bytes_0_t62 = 64'b0000000000000000000000000000000000000000000000000000000000000100;
    FSM_sub_bytes_0_t63 = FSM_sub_bytes_0_t62[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t64 = 64'b0000000000000000000000000000000000000000000000000000000000000100;
    FSM_sub_bytes_0_t65 = FSM_sub_bytes_0_t64[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t66 = FSM_sub_bytes_0_t61[FSM_sub_bytes_0_t65 * 64 +: 64];
    FSM_sub_bytes_0_t67 = FSM_sub_bytes_0_t66[6'b0 * 1 +: 8 * 1];
    FSM_sub_bytes_0_t68 = FSM_sub_bytes_0_t31[FSM_sub_bytes_0_t67 * 64 +: 64];
    FSM_sub_bytes_0_t69 = FSM_sub_bytes_0_t61;
    FSM_sub_bytes_0_t69[FSM_sub_bytes_0_t63 * 64 +: 64] = FSM_sub_bytes_0_t68;
    FSM_sub_bytes_0_t70 = 64'b0000000000000000000000000000000000000000000000000000000000000101;
    FSM_sub_bytes_0_t71 = FSM_sub_bytes_0_t70[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t72 = 64'b0000000000000000000000000000000000000000000000000000000000000101;
    FSM_sub_bytes_0_t73 = FSM_sub_bytes_0_t72[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t74 = FSM_sub_bytes_0_t69[FSM_sub_bytes_0_t73 * 64 +: 64];
    FSM_sub_bytes_0_t75 = FSM_sub_bytes_0_t74[6'b0 * 1 +: 8 * 1];
    FSM_sub_bytes_0_t76 = FSM_sub_bytes_0_t31[FSM_sub_bytes_0_t75 * 64 +: 64];
    FSM_sub_bytes_0_t77 = FSM_sub_bytes_0_t69;
    FSM_sub_bytes_0_t77[FSM_sub_bytes_0_t71 * 64 +: 64] = FSM_sub_bytes_0_t76;
    FSM_sub_bytes_0_t78 = 64'b0000000000000000000000000000000000000000000000000000000000000110;
    FSM_sub_bytes_0_t79 = FSM_sub_bytes_0_t78[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t80 = 64'b0000000000000000000000000000000000000000000000000000000000000110;
    FSM_sub_bytes_0_t81 = FSM_sub_bytes_0_t80[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t82 = FSM_sub_bytes_0_t77[FSM_sub_bytes_0_t81 * 64 +: 64];
    FSM_sub_bytes_0_t83 = FSM_sub_bytes_0_t82[6'b0 * 1 +: 8 * 1];
    FSM_sub_bytes_0_t84 = FSM_sub_bytes_0_t31[FSM_sub_bytes_0_t83 * 64 +: 64];
    FSM_sub_bytes_0_t85 = FSM_sub_bytes_0_t77;
    FSM_sub_bytes_0_t85[FSM_sub_bytes_0_t79 * 64 +: 64] = FSM_sub_bytes_0_t84;
    FSM_sub_bytes_0_t86 = 64'b0000000000000000000000000000000000000000000000000000000000000111;
    FSM_sub_bytes_0_t87 = FSM_sub_bytes_0_t86[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t88 = 64'b0000000000000000000000000000000000000000000000000000000000000111;
    FSM_sub_bytes_0_t89 = FSM_sub_bytes_0_t88[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t90 = FSM_sub_bytes_0_t85[FSM_sub_bytes_0_t89 * 64 +: 64];
    FSM_sub_bytes_0_t91 = FSM_sub_bytes_0_t90[6'b0 * 1 +: 8 * 1];
    FSM_sub_bytes_0_t92 = FSM_sub_bytes_0_t31[FSM_sub_bytes_0_t91 * 64 +: 64];
    FSM_sub_bytes_0_t93 = FSM_sub_bytes_0_t85;
    FSM_sub_bytes_0_t93[FSM_sub_bytes_0_t87 * 64 +: 64] = FSM_sub_bytes_0_t92;
    FSM_sub_bytes_0_t94 = 64'b0000000000000000000000000000000000000000000000000000000000001000;
    FSM_sub_bytes_0_t95 = FSM_sub_bytes_0_t94[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t96 = 64'b0000000000000000000000000000000000000000000000000000000000001000;
    FSM_sub_bytes_0_t97 = FSM_sub_bytes_0_t96[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t98 = FSM_sub_bytes_0_t93[FSM_sub_bytes_0_t97 * 64 +: 64];
    FSM_sub_bytes_0_t99 = FSM_sub_bytes_0_t98[6'b0 * 1 +: 8 * 1];
    FSM_sub_bytes_0_t100 = FSM_sub_bytes_0_t31[FSM_sub_bytes_0_t99 * 64 +: 64];
    FSM_sub_bytes_0_t101 = FSM_sub_bytes_0_t93;
    FSM_sub_bytes_0_t101[FSM_sub_bytes_0_t95 * 64 +: 64] = FSM_sub_bytes_0_t100;
    FSM_sub_bytes_0_t102 = 64'b0000000000000000000000000000000000000000000000000000000000001001;
    FSM_sub_bytes_0_t103 = FSM_sub_bytes_0_t102[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t104 = 64'b0000000000000000000000000000000000000000000000000000000000001001;
    FSM_sub_bytes_0_t105 = FSM_sub_bytes_0_t104[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t106 = FSM_sub_bytes_0_t101[FSM_sub_bytes_0_t105 * 64 +: 64];
    FSM_sub_bytes_0_t107 = FSM_sub_bytes_0_t106[6'b0 * 1 +: 8 * 1];
    FSM_sub_bytes_0_t108 = FSM_sub_bytes_0_t31[FSM_sub_bytes_0_t107 * 64 +: 64];
    FSM_sub_bytes_0_t109 = FSM_sub_bytes_0_t101;
    FSM_sub_bytes_0_t109[FSM_sub_bytes_0_t103 * 64 +: 64] = FSM_sub_bytes_0_t108;
    FSM_sub_bytes_0_t110 = 64'b0000000000000000000000000000000000000000000000000000000000001010;
    FSM_sub_bytes_0_t111 = FSM_sub_bytes_0_t110[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t112 = 64'b0000000000000000000000000000000000000000000000000000000000001010;
    FSM_sub_bytes_0_t113 = FSM_sub_bytes_0_t112[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t114 = FSM_sub_bytes_0_t109[FSM_sub_bytes_0_t113 * 64 +: 64];
    FSM_sub_bytes_0_t115 = FSM_sub_bytes_0_t114[6'b0 * 1 +: 8 * 1];
    FSM_sub_bytes_0_t116 = FSM_sub_bytes_0_t31[FSM_sub_bytes_0_t115 * 64 +: 64];
    FSM_sub_bytes_0_t117 = FSM_sub_bytes_0_t109;
    FSM_sub_bytes_0_t117[FSM_sub_bytes_0_t111 * 64 +: 64] = FSM_sub_bytes_0_t116;
    FSM_sub_bytes_0_t118 = 64'b0000000000000000000000000000000000000000000000000000000000001011;
    FSM_sub_bytes_0_t119 = FSM_sub_bytes_0_t118[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t120 = 64'b0000000000000000000000000000000000000000000000000000000000001011;
    FSM_sub_bytes_0_t121 = FSM_sub_bytes_0_t120[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t122 = FSM_sub_bytes_0_t117[FSM_sub_bytes_0_t121 * 64 +: 64];
    FSM_sub_bytes_0_t123 = FSM_sub_bytes_0_t122[6'b0 * 1 +: 8 * 1];
    FSM_sub_bytes_0_t124 = FSM_sub_bytes_0_t31[FSM_sub_bytes_0_t123 * 64 +: 64];
    FSM_sub_bytes_0_t125 = FSM_sub_bytes_0_t117;
    FSM_sub_bytes_0_t125[FSM_sub_bytes_0_t119 * 64 +: 64] = FSM_sub_bytes_0_t124;
    FSM_sub_bytes_0_t126 = 64'b0000000000000000000000000000000000000000000000000000000000001100;
    FSM_sub_bytes_0_t127 = FSM_sub_bytes_0_t126[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t128 = 64'b0000000000000000000000000000000000000000000000000000000000001100;
    FSM_sub_bytes_0_t129 = FSM_sub_bytes_0_t128[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t130 = FSM_sub_bytes_0_t125[FSM_sub_bytes_0_t129 * 64 +: 64];
    FSM_sub_bytes_0_t131 = FSM_sub_bytes_0_t130[6'b0 * 1 +: 8 * 1];
    FSM_sub_bytes_0_t132 = FSM_sub_bytes_0_t31[FSM_sub_bytes_0_t131 * 64 +: 64];
    FSM_sub_bytes_0_t133 = FSM_sub_bytes_0_t125;
    FSM_sub_bytes_0_t133[FSM_sub_bytes_0_t127 * 64 +: 64] = FSM_sub_bytes_0_t132;
    FSM_sub_bytes_0_t134 = 64'b0000000000000000000000000000000000000000000000000000000000001101;
    FSM_sub_bytes_0_t135 = FSM_sub_bytes_0_t134[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t136 = 64'b0000000000000000000000000000000000000000000000000000000000001101;
    FSM_sub_bytes_0_t137 = FSM_sub_bytes_0_t136[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t138 = FSM_sub_bytes_0_t133[FSM_sub_bytes_0_t137 * 64 +: 64];
    FSM_sub_bytes_0_t139 = FSM_sub_bytes_0_t138[6'b0 * 1 +: 8 * 1];
    FSM_sub_bytes_0_t140 = FSM_sub_bytes_0_t31[FSM_sub_bytes_0_t139 * 64 +: 64];
    FSM_sub_bytes_0_t141 = FSM_sub_bytes_0_t133;
    FSM_sub_bytes_0_t141[FSM_sub_bytes_0_t135 * 64 +: 64] = FSM_sub_bytes_0_t140;
    FSM_sub_bytes_0_t142 = 64'b0000000000000000000000000000000000000000000000000000000000001110;
    FSM_sub_bytes_0_t143 = FSM_sub_bytes_0_t142[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t144 = 64'b0000000000000000000000000000000000000000000000000000000000001110;
    FSM_sub_bytes_0_t145 = FSM_sub_bytes_0_t144[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t146 = FSM_sub_bytes_0_t141[FSM_sub_bytes_0_t145 * 64 +: 64];
    FSM_sub_bytes_0_t147 = FSM_sub_bytes_0_t146[6'b0 * 1 +: 8 * 1];
    FSM_sub_bytes_0_t148 = FSM_sub_bytes_0_t31[FSM_sub_bytes_0_t147 * 64 +: 64];
    FSM_sub_bytes_0_t149 = FSM_sub_bytes_0_t141;
    FSM_sub_bytes_0_t149[FSM_sub_bytes_0_t143 * 64 +: 64] = FSM_sub_bytes_0_t148;
    FSM_sub_bytes_0_t150 = 64'b0000000000000000000000000000000000000000000000000000000000001111;
    FSM_sub_bytes_0_t151 = FSM_sub_bytes_0_t150[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t152 = 64'b0000000000000000000000000000000000000000000000000000000000001111;
    FSM_sub_bytes_0_t153 = FSM_sub_bytes_0_t152[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t154 = FSM_sub_bytes_0_t149[FSM_sub_bytes_0_t153 * 64 +: 64];
    FSM_sub_bytes_0_t155 = FSM_sub_bytes_0_t154[6'b0 * 1 +: 8 * 1];
    FSM_sub_bytes_0_t156 = FSM_sub_bytes_0_t31[FSM_sub_bytes_0_t155 * 64 +: 64];
    FSM_sub_bytes_0_t157 = FSM_sub_bytes_0_t149;
    FSM_sub_bytes_0_t157[FSM_sub_bytes_0_t151 * 64 +: 64] = FSM_sub_bytes_0_t156;
    FSM_sub_bytes_0_t158 = 64'b0;
    FSM_sub_bytes_0_t159 = FSM_sub_bytes_0_t158[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t160 = FSM_sub_bytes_0_t157[FSM_sub_bytes_0_t159 * 64 +: 64];
    FSM_sub_bytes_0_t161 = 64'b0000000000000000000000000000000000000000000000000000000000000001;
    FSM_sub_bytes_0_t162 = FSM_sub_bytes_0_t161[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t163 = FSM_sub_bytes_0_t157[FSM_sub_bytes_0_t162 * 64 +: 64];
    FSM_sub_bytes_0_t164 = 64'b0000000000000000000000000000000000000000000000000000000000001000;
    FSM_sub_bytes_0_t165 = FSM_sub_bytes_0_t164[6'b0 * 1 +: 6 * 1];
    FSM_sub_bytes_0_t166 = 64'b0000000000000000000000000000000000000000000000000000000000000010;
    FSM_sub_bytes_0_t167 = FSM_sub_bytes_0_t166[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t168 = FSM_sub_bytes_0_t157[FSM_sub_bytes_0_t167 * 64 +: 64];
    FSM_sub_bytes_0_t169 = 64'b0000000000000000000000000000000000000000000000000000000000010000;
    FSM_sub_bytes_0_t170 = FSM_sub_bytes_0_t169[6'b0 * 1 +: 6 * 1];
    FSM_sub_bytes_0_t171 = 64'b0000000000000000000000000000000000000000000000000000000000000011;
    FSM_sub_bytes_0_t172 = FSM_sub_bytes_0_t171[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t173 = FSM_sub_bytes_0_t157[FSM_sub_bytes_0_t172 * 64 +: 64];
    FSM_sub_bytes_0_t174 = 64'b0000000000000000000000000000000000000000000000000000000000011000;
    FSM_sub_bytes_0_t175 = FSM_sub_bytes_0_t174[6'b0 * 1 +: 6 * 1];
    FSM_sub_bytes_0_t176 = 64'b0000000000000000000000000000000000000000000000000000000000000100;
    FSM_sub_bytes_0_t177 = FSM_sub_bytes_0_t176[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t178 = FSM_sub_bytes_0_t157[FSM_sub_bytes_0_t177 * 64 +: 64];
    FSM_sub_bytes_0_t179 = 64'b0000000000000000000000000000000000000000000000000000000000100000;
    FSM_sub_bytes_0_t180 = FSM_sub_bytes_0_t179[6'b0 * 1 +: 6 * 1];
    FSM_sub_bytes_0_t181 = 64'b0000000000000000000000000000000000000000000000000000000000000101;
    FSM_sub_bytes_0_t182 = FSM_sub_bytes_0_t181[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t183 = FSM_sub_bytes_0_t157[FSM_sub_bytes_0_t182 * 64 +: 64];
    FSM_sub_bytes_0_t184 = 64'b0000000000000000000000000000000000000000000000000000000000101000;
    FSM_sub_bytes_0_t185 = FSM_sub_bytes_0_t184[6'b0 * 1 +: 6 * 1];
    FSM_sub_bytes_0_t186 = 64'b0000000000000000000000000000000000000000000000000000000000000110;
    FSM_sub_bytes_0_t187 = FSM_sub_bytes_0_t186[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t188 = FSM_sub_bytes_0_t157[FSM_sub_bytes_0_t187 * 64 +: 64];
    FSM_sub_bytes_0_t189 = 64'b0000000000000000000000000000000000000000000000000000000000110000;
    FSM_sub_bytes_0_t190 = FSM_sub_bytes_0_t189[6'b0 * 1 +: 6 * 1];
    FSM_sub_bytes_0_t191 = 64'b0000000000000000000000000000000000000000000000000000000000000111;
    FSM_sub_bytes_0_t192 = FSM_sub_bytes_0_t191[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t193 = FSM_sub_bytes_0_t157[FSM_sub_bytes_0_t192 * 64 +: 64];
    FSM_sub_bytes_0_t194 = 64'b0000000000000000000000000000000000000000000000000000000000111000;
    FSM_sub_bytes_0_t195 = FSM_sub_bytes_0_t194[6'b0 * 1 +: 6 * 1];
    FSM_sub_bytes_0_t196 = 64'b0000000000000000000000000000000000000000000000000000000000001000;
    FSM_sub_bytes_0_t197 = FSM_sub_bytes_0_t196[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t198 = FSM_sub_bytes_0_t157[FSM_sub_bytes_0_t197 * 64 +: 64];
    FSM_sub_bytes_0_t199 = 64'b0000000000000000000000000000000000000000000000000000000000001001;
    FSM_sub_bytes_0_t200 = FSM_sub_bytes_0_t199[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t201 = FSM_sub_bytes_0_t157[FSM_sub_bytes_0_t200 * 64 +: 64];
    FSM_sub_bytes_0_t202 = 64'b0000000000000000000000000000000000000000000000000000000000001000;
    FSM_sub_bytes_0_t203 = FSM_sub_bytes_0_t202[6'b0 * 1 +: 6 * 1];
    FSM_sub_bytes_0_t204 = 64'b0000000000000000000000000000000000000000000000000000000000001010;
    FSM_sub_bytes_0_t205 = FSM_sub_bytes_0_t204[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t206 = FSM_sub_bytes_0_t157[FSM_sub_bytes_0_t205 * 64 +: 64];
    FSM_sub_bytes_0_t207 = 64'b0000000000000000000000000000000000000000000000000000000000010000;
    FSM_sub_bytes_0_t208 = FSM_sub_bytes_0_t207[6'b0 * 1 +: 6 * 1];
    FSM_sub_bytes_0_t209 = 64'b0000000000000000000000000000000000000000000000000000000000001011;
    FSM_sub_bytes_0_t210 = FSM_sub_bytes_0_t209[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t211 = FSM_sub_bytes_0_t157[FSM_sub_bytes_0_t210 * 64 +: 64];
    FSM_sub_bytes_0_t212 = 64'b0000000000000000000000000000000000000000000000000000000000011000;
    FSM_sub_bytes_0_t213 = FSM_sub_bytes_0_t212[6'b0 * 1 +: 6 * 1];
    FSM_sub_bytes_0_t214 = 64'b0000000000000000000000000000000000000000000000000000000000001100;
    FSM_sub_bytes_0_t215 = FSM_sub_bytes_0_t214[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t216 = FSM_sub_bytes_0_t157[FSM_sub_bytes_0_t215 * 64 +: 64];
    FSM_sub_bytes_0_t217 = 64'b0000000000000000000000000000000000000000000000000000000000100000;
    FSM_sub_bytes_0_t218 = FSM_sub_bytes_0_t217[6'b0 * 1 +: 6 * 1];
    FSM_sub_bytes_0_t219 = 64'b0000000000000000000000000000000000000000000000000000000000001101;
    FSM_sub_bytes_0_t220 = FSM_sub_bytes_0_t219[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t221 = FSM_sub_bytes_0_t157[FSM_sub_bytes_0_t220 * 64 +: 64];
    FSM_sub_bytes_0_t222 = 64'b0000000000000000000000000000000000000000000000000000000000101000;
    FSM_sub_bytes_0_t223 = FSM_sub_bytes_0_t222[6'b0 * 1 +: 6 * 1];
    FSM_sub_bytes_0_t224 = 64'b0000000000000000000000000000000000000000000000000000000000001110;
    FSM_sub_bytes_0_t225 = FSM_sub_bytes_0_t224[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t226 = FSM_sub_bytes_0_t157[FSM_sub_bytes_0_t225 * 64 +: 64];
    FSM_sub_bytes_0_t227 = 64'b0000000000000000000000000000000000000000000000000000000000110000;
    FSM_sub_bytes_0_t228 = FSM_sub_bytes_0_t227[6'b0 * 1 +: 6 * 1];
    FSM_sub_bytes_0_t229 = 64'b0000000000000000000000000000000000000000000000000000000000001111;
    FSM_sub_bytes_0_t230 = FSM_sub_bytes_0_t229[6'b0 * 1 +: 4 * 1];
    FSM_sub_bytes_0_t231 = FSM_sub_bytes_0_t157[FSM_sub_bytes_0_t230 * 64 +: 64];
    FSM_sub_bytes_0_t232 = 64'b0000000000000000000000000000000000000000000000000000000000111000;
    FSM_sub_bytes_0_t233 = FSM_sub_bytes_0_t232[6'b0 * 1 +: 6 * 1];
end

assign FSM_sub_bytes_0_in_ready = 1'b1;

always @(posedge clk) begin
    FSM_sub_bytes_0_st_dummy_reg <= FSM_sub_bytes_0_st_dummy_reg;
    if (rst) begin
        FSM_sub_bytes_0_st_dummy_reg <= 64'b0;
    end
end
/* End submodules of sub_bytes */
/* End module sub_bytes */
endgenerate
endmodule
