package acc_pkg;
	typedef struct packed {
		logic dummy;
	} acc_config_t;
endpackage : acc_pkg