`timescale 1ns / 1ps

module dct_8x8_stage_8_inner
(
    input wire clk,
    input wire rst,
    input wire [2048-1:0] i_data_in,
    input wire i_valid,
    output wire i_ready,
    output wire [2048-1:0] o_data_out,
    output wire o_valid,
    input wire o_ready
);

generate
/*
    Begin module dct_8x8_stage_8
*/
/*
    Wires declared by dct_8x8_stage_8
*/
wire FSM_dct_8x8_stage_8_0_in_ready;
wire FSM_dct_8x8_stage_8_0_out_valid;
/* End wires declared by dct_8x8_stage_8 */

/*
    Submodules of dct_8x8_stage_8
*/
reg [32-1:0] FSM_dct_8x8_stage_8_0_st_dummy_reg = 32'b0;

reg [32-1:0] FSM_dct_8x8_stage_8_0_t0;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t1;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t2;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t3;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t4;
reg [2048-1:0] FSM_dct_8x8_stage_8_0_t5;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t6;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t7;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t8;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t9;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t10;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t11;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t12;
reg [2048-1:0] FSM_dct_8x8_stage_8_0_t13;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t14;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t15;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t16;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t17;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t18;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t19;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t20;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t21;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t22;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t23;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t24;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t25;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t26;
reg [2048-1:0] FSM_dct_8x8_stage_8_0_t27;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t28;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t29;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t30;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t31;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t32;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t33;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t34;
reg [2048-1:0] FSM_dct_8x8_stage_8_0_t35;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t36;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t37;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t38;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t39;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t40;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t41;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t42;
reg [2048-1:0] FSM_dct_8x8_stage_8_0_t43;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t44;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t45;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t46;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t47;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t48;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t49;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t50;
reg [2048-1:0] FSM_dct_8x8_stage_8_0_t51;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t52;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t53;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t54;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t55;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t56;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t57;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t58;
reg [2048-1:0] FSM_dct_8x8_stage_8_0_t59;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t60;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t61;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t62;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t63;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t64;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t65;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t66;
reg [2048-1:0] FSM_dct_8x8_stage_8_0_t67;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t68;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t69;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t70;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t71;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t72;
reg [2048-1:0] FSM_dct_8x8_stage_8_0_t73;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t74;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t75;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t76;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t77;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t78;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t79;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t80;
reg [2048-1:0] FSM_dct_8x8_stage_8_0_t81;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t82;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t83;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t84;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t85;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t86;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t87;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t88;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t89;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t90;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t91;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t92;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t93;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t94;
reg [2048-1:0] FSM_dct_8x8_stage_8_0_t95;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t96;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t97;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t98;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t99;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t100;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t101;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t102;
reg [2048-1:0] FSM_dct_8x8_stage_8_0_t103;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t104;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t105;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t106;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t107;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t108;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t109;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t110;
reg [2048-1:0] FSM_dct_8x8_stage_8_0_t111;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t112;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t113;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t114;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t115;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t116;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t117;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t118;
reg [2048-1:0] FSM_dct_8x8_stage_8_0_t119;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t120;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t121;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t122;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t123;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t124;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t125;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t126;
reg [2048-1:0] FSM_dct_8x8_stage_8_0_t127;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t128;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t129;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t130;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t131;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t132;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t133;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t134;
reg [2048-1:0] FSM_dct_8x8_stage_8_0_t135;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t136;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t137;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t138;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t139;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t140;
reg [2048-1:0] FSM_dct_8x8_stage_8_0_t141;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t142;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t143;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t144;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t145;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t146;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t147;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t148;
reg [2048-1:0] FSM_dct_8x8_stage_8_0_t149;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t150;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t151;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t152;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t153;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t154;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t155;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t156;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t157;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t158;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t159;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t160;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t161;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t162;
reg [2048-1:0] FSM_dct_8x8_stage_8_0_t163;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t164;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t165;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t166;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t167;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t168;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t169;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t170;
reg [2048-1:0] FSM_dct_8x8_stage_8_0_t171;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t172;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t173;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t174;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t175;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t176;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t177;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t178;
reg [2048-1:0] FSM_dct_8x8_stage_8_0_t179;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t180;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t181;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t182;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t183;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t184;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t185;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t186;
reg [2048-1:0] FSM_dct_8x8_stage_8_0_t187;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t188;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t189;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t190;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t191;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t192;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t193;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t194;
reg [2048-1:0] FSM_dct_8x8_stage_8_0_t195;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t196;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t197;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t198;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t199;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t200;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t201;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t202;
reg [2048-1:0] FSM_dct_8x8_stage_8_0_t203;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t204;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t205;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t206;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t207;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t208;
reg [2048-1:0] FSM_dct_8x8_stage_8_0_t209;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t210;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t211;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t212;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t213;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t214;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t215;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t216;
reg [2048-1:0] FSM_dct_8x8_stage_8_0_t217;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t218;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t219;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t220;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t221;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t222;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t223;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t224;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t225;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t226;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t227;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t228;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t229;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t230;
reg [2048-1:0] FSM_dct_8x8_stage_8_0_t231;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t232;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t233;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t234;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t235;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t236;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t237;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t238;
reg [2048-1:0] FSM_dct_8x8_stage_8_0_t239;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t240;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t241;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t242;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t243;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t244;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t245;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t246;
reg [2048-1:0] FSM_dct_8x8_stage_8_0_t247;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t248;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t249;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t250;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t251;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t252;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t253;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t254;
reg [2048-1:0] FSM_dct_8x8_stage_8_0_t255;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t256;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t257;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t258;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t259;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t260;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t261;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t262;
reg [2048-1:0] FSM_dct_8x8_stage_8_0_t263;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t264;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t265;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t266;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t267;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t268;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t269;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t270;
reg [2048-1:0] FSM_dct_8x8_stage_8_0_t271;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t272;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t273;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t274;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t275;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t276;
reg [2048-1:0] FSM_dct_8x8_stage_8_0_t277;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t278;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t279;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t280;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t281;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t282;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t283;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t284;
reg [2048-1:0] FSM_dct_8x8_stage_8_0_t285;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t286;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t287;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t288;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t289;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t290;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t291;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t292;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t293;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t294;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t295;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t296;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t297;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t298;
reg [2048-1:0] FSM_dct_8x8_stage_8_0_t299;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t300;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t301;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t302;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t303;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t304;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t305;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t306;
reg [2048-1:0] FSM_dct_8x8_stage_8_0_t307;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t308;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t309;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t310;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t311;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t312;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t313;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t314;
reg [2048-1:0] FSM_dct_8x8_stage_8_0_t315;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t316;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t317;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t318;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t319;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t320;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t321;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t322;
reg [2048-1:0] FSM_dct_8x8_stage_8_0_t323;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t324;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t325;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t326;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t327;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t328;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t329;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t330;
reg [2048-1:0] FSM_dct_8x8_stage_8_0_t331;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t332;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t333;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t334;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t335;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t336;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t337;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t338;
reg [2048-1:0] FSM_dct_8x8_stage_8_0_t339;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t340;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t341;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t342;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t343;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t344;
reg [2048-1:0] FSM_dct_8x8_stage_8_0_t345;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t346;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t347;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t348;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t349;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t350;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t351;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t352;
reg [2048-1:0] FSM_dct_8x8_stage_8_0_t353;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t354;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t355;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t356;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t357;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t358;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t359;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t360;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t361;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t362;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t363;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t364;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t365;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t366;
reg [2048-1:0] FSM_dct_8x8_stage_8_0_t367;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t368;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t369;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t370;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t371;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t372;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t373;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t374;
reg [2048-1:0] FSM_dct_8x8_stage_8_0_t375;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t376;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t377;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t378;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t379;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t380;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t381;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t382;
reg [2048-1:0] FSM_dct_8x8_stage_8_0_t383;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t384;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t385;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t386;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t387;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t388;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t389;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t390;
reg [2048-1:0] FSM_dct_8x8_stage_8_0_t391;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t392;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t393;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t394;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t395;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t396;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t397;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t398;
reg [2048-1:0] FSM_dct_8x8_stage_8_0_t399;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t400;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t401;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t402;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t403;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t404;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t405;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t406;
reg [2048-1:0] FSM_dct_8x8_stage_8_0_t407;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t408;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t409;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t410;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t411;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t412;
reg [2048-1:0] FSM_dct_8x8_stage_8_0_t413;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t414;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t415;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t416;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t417;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t418;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t419;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t420;
reg [2048-1:0] FSM_dct_8x8_stage_8_0_t421;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t422;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t423;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t424;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t425;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t426;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t427;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t428;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t429;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t430;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t431;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t432;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t433;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t434;
reg [2048-1:0] FSM_dct_8x8_stage_8_0_t435;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t436;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t437;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t438;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t439;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t440;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t441;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t442;
reg [2048-1:0] FSM_dct_8x8_stage_8_0_t443;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t444;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t445;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t446;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t447;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t448;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t449;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t450;
reg [2048-1:0] FSM_dct_8x8_stage_8_0_t451;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t452;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t453;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t454;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t455;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t456;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t457;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t458;
reg [2048-1:0] FSM_dct_8x8_stage_8_0_t459;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t460;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t461;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t462;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t463;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t464;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t465;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t466;
reg [2048-1:0] FSM_dct_8x8_stage_8_0_t467;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t468;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t469;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t470;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t471;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t472;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t473;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t474;
reg [2048-1:0] FSM_dct_8x8_stage_8_0_t475;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t476;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t477;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t478;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t479;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t480;
reg [2048-1:0] FSM_dct_8x8_stage_8_0_t481;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t482;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t483;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t484;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t485;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t486;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t487;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t488;
reg [2048-1:0] FSM_dct_8x8_stage_8_0_t489;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t490;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t491;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t492;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t493;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t494;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t495;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t496;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t497;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t498;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t499;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t500;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t501;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t502;
reg [2048-1:0] FSM_dct_8x8_stage_8_0_t503;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t504;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t505;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t506;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t507;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t508;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t509;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t510;
reg [2048-1:0] FSM_dct_8x8_stage_8_0_t511;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t512;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t513;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t514;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t515;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t516;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t517;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t518;
reg [2048-1:0] FSM_dct_8x8_stage_8_0_t519;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t520;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t521;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t522;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t523;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t524;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t525;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t526;
reg [2048-1:0] FSM_dct_8x8_stage_8_0_t527;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t528;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t529;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t530;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t531;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t532;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t533;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t534;
reg [2048-1:0] FSM_dct_8x8_stage_8_0_t535;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t536;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t537;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t538;
reg [33-1:0] FSM_dct_8x8_stage_8_0_t539;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t540;
reg [6-1:0] FSM_dct_8x8_stage_8_0_t541;
reg [32-1:0] FSM_dct_8x8_stage_8_0_t542;
reg [2048-1:0] FSM_dct_8x8_stage_8_0_t543;

/*
    Wiring by dct_8x8_stage_8
*/
assign i_ready = FSM_dct_8x8_stage_8_0_in_ready;
assign o_data_out = FSM_dct_8x8_stage_8_0_t543;
assign o_valid = FSM_dct_8x8_stage_8_0_out_valid;
/* End wiring by dct_8x8_stage_8 */

assign FSM_dct_8x8_stage_8_0_out_valid = 1'b1;

initial begin
    FSM_dct_8x8_stage_8_0_t0 = 32'b0;
    FSM_dct_8x8_stage_8_0_t1 = FSM_dct_8x8_stage_8_0_t0[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t2 = 32'b0;
    FSM_dct_8x8_stage_8_0_t3 = FSM_dct_8x8_stage_8_0_t2[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t4 = i_data_in[FSM_dct_8x8_stage_8_0_t3 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t5 = 2048'b0;
    FSM_dct_8x8_stage_8_0_t5[FSM_dct_8x8_stage_8_0_t1 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t4;
    FSM_dct_8x8_stage_8_0_t6 = 32'b00000000000000000000000000001000 + 32'b0;
    FSM_dct_8x8_stage_8_0_t7 = FSM_dct_8x8_stage_8_0_t6[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t8 = FSM_dct_8x8_stage_8_0_t7[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t9 = 32'b00000000000000000000000000001000 + 32'b0;
    FSM_dct_8x8_stage_8_0_t10 = FSM_dct_8x8_stage_8_0_t9[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t11 = FSM_dct_8x8_stage_8_0_t10[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t12 = i_data_in[FSM_dct_8x8_stage_8_0_t11 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t13 = FSM_dct_8x8_stage_8_0_t5;
    FSM_dct_8x8_stage_8_0_t13[FSM_dct_8x8_stage_8_0_t8 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t12;
    FSM_dct_8x8_stage_8_0_t14 = 32'b00000000000000000000000000010000 + 32'b0;
    FSM_dct_8x8_stage_8_0_t15 = FSM_dct_8x8_stage_8_0_t14[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t16 = FSM_dct_8x8_stage_8_0_t15[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t17 = 32'b00000000000000000000000000010000 + 32'b0;
    FSM_dct_8x8_stage_8_0_t18 = FSM_dct_8x8_stage_8_0_t17[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t19 = FSM_dct_8x8_stage_8_0_t18[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t20 = i_data_in[FSM_dct_8x8_stage_8_0_t19 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t21 = 32'b00000000000000000000000000011000 + 32'b0;
    FSM_dct_8x8_stage_8_0_t22 = FSM_dct_8x8_stage_8_0_t21[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t23 = FSM_dct_8x8_stage_8_0_t22[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t24 = i_data_in[FSM_dct_8x8_stage_8_0_t23 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t25 = FSM_dct_8x8_stage_8_0_t20 + FSM_dct_8x8_stage_8_0_t24;
    FSM_dct_8x8_stage_8_0_t26 = FSM_dct_8x8_stage_8_0_t25[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t27 = FSM_dct_8x8_stage_8_0_t13;
    FSM_dct_8x8_stage_8_0_t27[FSM_dct_8x8_stage_8_0_t16 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t26;
    FSM_dct_8x8_stage_8_0_t28 = 32'b00000000000000000000000000011000 + 32'b0;
    FSM_dct_8x8_stage_8_0_t29 = FSM_dct_8x8_stage_8_0_t28[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t30 = FSM_dct_8x8_stage_8_0_t29[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t31 = 32'b00000000000000000000000000011000 + 32'b0;
    FSM_dct_8x8_stage_8_0_t32 = FSM_dct_8x8_stage_8_0_t31[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t33 = FSM_dct_8x8_stage_8_0_t32[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t34 = i_data_in[FSM_dct_8x8_stage_8_0_t33 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t35 = FSM_dct_8x8_stage_8_0_t27;
    FSM_dct_8x8_stage_8_0_t35[FSM_dct_8x8_stage_8_0_t30 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t34;
    FSM_dct_8x8_stage_8_0_t36 = 32'b00000000000000000000000000100000 + 32'b0;
    FSM_dct_8x8_stage_8_0_t37 = FSM_dct_8x8_stage_8_0_t36[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t38 = FSM_dct_8x8_stage_8_0_t37[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t39 = 32'b00000000000000000000000000100000 + 32'b0;
    FSM_dct_8x8_stage_8_0_t40 = FSM_dct_8x8_stage_8_0_t39[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t41 = FSM_dct_8x8_stage_8_0_t40[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t42 = i_data_in[FSM_dct_8x8_stage_8_0_t41 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t43 = FSM_dct_8x8_stage_8_0_t35;
    FSM_dct_8x8_stage_8_0_t43[FSM_dct_8x8_stage_8_0_t38 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t42;
    FSM_dct_8x8_stage_8_0_t44 = 32'b00000000000000000000000000101000 + 32'b0;
    FSM_dct_8x8_stage_8_0_t45 = FSM_dct_8x8_stage_8_0_t44[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t46 = FSM_dct_8x8_stage_8_0_t45[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t47 = 32'b00000000000000000000000000101000 + 32'b0;
    FSM_dct_8x8_stage_8_0_t48 = FSM_dct_8x8_stage_8_0_t47[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t49 = FSM_dct_8x8_stage_8_0_t48[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t50 = i_data_in[FSM_dct_8x8_stage_8_0_t49 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t51 = FSM_dct_8x8_stage_8_0_t43;
    FSM_dct_8x8_stage_8_0_t51[FSM_dct_8x8_stage_8_0_t46 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t50;
    FSM_dct_8x8_stage_8_0_t52 = 32'b00000000000000000000000000110000 + 32'b0;
    FSM_dct_8x8_stage_8_0_t53 = FSM_dct_8x8_stage_8_0_t52[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t54 = FSM_dct_8x8_stage_8_0_t53[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t55 = 32'b00000000000000000000000000110000 + 32'b0;
    FSM_dct_8x8_stage_8_0_t56 = FSM_dct_8x8_stage_8_0_t55[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t57 = FSM_dct_8x8_stage_8_0_t56[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t58 = i_data_in[FSM_dct_8x8_stage_8_0_t57 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t59 = FSM_dct_8x8_stage_8_0_t51;
    FSM_dct_8x8_stage_8_0_t59[FSM_dct_8x8_stage_8_0_t54 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t58;
    FSM_dct_8x8_stage_8_0_t60 = 32'b00000000000000000000000000111000 + 32'b0;
    FSM_dct_8x8_stage_8_0_t61 = FSM_dct_8x8_stage_8_0_t60[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t62 = FSM_dct_8x8_stage_8_0_t61[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t63 = 32'b00000000000000000000000000111000 + 32'b0;
    FSM_dct_8x8_stage_8_0_t64 = FSM_dct_8x8_stage_8_0_t63[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t65 = FSM_dct_8x8_stage_8_0_t64[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t66 = i_data_in[FSM_dct_8x8_stage_8_0_t65 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t67 = FSM_dct_8x8_stage_8_0_t59;
    FSM_dct_8x8_stage_8_0_t67[FSM_dct_8x8_stage_8_0_t62 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t66;
    FSM_dct_8x8_stage_8_0_t68 = 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_8_0_t69 = FSM_dct_8x8_stage_8_0_t68[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t70 = 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_8_0_t71 = FSM_dct_8x8_stage_8_0_t70[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t72 = i_data_in[FSM_dct_8x8_stage_8_0_t71 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t73 = FSM_dct_8x8_stage_8_0_t67;
    FSM_dct_8x8_stage_8_0_t73[FSM_dct_8x8_stage_8_0_t69 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t72;
    FSM_dct_8x8_stage_8_0_t74 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_8_0_t75 = FSM_dct_8x8_stage_8_0_t74[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t76 = FSM_dct_8x8_stage_8_0_t75[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t77 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_8_0_t78 = FSM_dct_8x8_stage_8_0_t77[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t79 = FSM_dct_8x8_stage_8_0_t78[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t80 = i_data_in[FSM_dct_8x8_stage_8_0_t79 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t81 = FSM_dct_8x8_stage_8_0_t73;
    FSM_dct_8x8_stage_8_0_t81[FSM_dct_8x8_stage_8_0_t76 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t80;
    FSM_dct_8x8_stage_8_0_t82 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_8_0_t83 = FSM_dct_8x8_stage_8_0_t82[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t84 = FSM_dct_8x8_stage_8_0_t83[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t85 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_8_0_t86 = FSM_dct_8x8_stage_8_0_t85[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t87 = FSM_dct_8x8_stage_8_0_t86[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t88 = i_data_in[FSM_dct_8x8_stage_8_0_t87 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t89 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_8_0_t90 = FSM_dct_8x8_stage_8_0_t89[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t91 = FSM_dct_8x8_stage_8_0_t90[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t92 = i_data_in[FSM_dct_8x8_stage_8_0_t91 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t93 = FSM_dct_8x8_stage_8_0_t88 + FSM_dct_8x8_stage_8_0_t92;
    FSM_dct_8x8_stage_8_0_t94 = FSM_dct_8x8_stage_8_0_t93[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t95 = FSM_dct_8x8_stage_8_0_t81;
    FSM_dct_8x8_stage_8_0_t95[FSM_dct_8x8_stage_8_0_t84 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t94;
    FSM_dct_8x8_stage_8_0_t96 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_8_0_t97 = FSM_dct_8x8_stage_8_0_t96[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t98 = FSM_dct_8x8_stage_8_0_t97[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t99 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_8_0_t100 = FSM_dct_8x8_stage_8_0_t99[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t101 = FSM_dct_8x8_stage_8_0_t100[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t102 = i_data_in[FSM_dct_8x8_stage_8_0_t101 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t103 = FSM_dct_8x8_stage_8_0_t95;
    FSM_dct_8x8_stage_8_0_t103[FSM_dct_8x8_stage_8_0_t98 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t102;
    FSM_dct_8x8_stage_8_0_t104 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_8_0_t105 = FSM_dct_8x8_stage_8_0_t104[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t106 = FSM_dct_8x8_stage_8_0_t105[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t107 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_8_0_t108 = FSM_dct_8x8_stage_8_0_t107[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t109 = FSM_dct_8x8_stage_8_0_t108[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t110 = i_data_in[FSM_dct_8x8_stage_8_0_t109 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t111 = FSM_dct_8x8_stage_8_0_t103;
    FSM_dct_8x8_stage_8_0_t111[FSM_dct_8x8_stage_8_0_t106 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t110;
    FSM_dct_8x8_stage_8_0_t112 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_8_0_t113 = FSM_dct_8x8_stage_8_0_t112[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t114 = FSM_dct_8x8_stage_8_0_t113[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t115 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_8_0_t116 = FSM_dct_8x8_stage_8_0_t115[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t117 = FSM_dct_8x8_stage_8_0_t116[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t118 = i_data_in[FSM_dct_8x8_stage_8_0_t117 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t119 = FSM_dct_8x8_stage_8_0_t111;
    FSM_dct_8x8_stage_8_0_t119[FSM_dct_8x8_stage_8_0_t114 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t118;
    FSM_dct_8x8_stage_8_0_t120 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_8_0_t121 = FSM_dct_8x8_stage_8_0_t120[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t122 = FSM_dct_8x8_stage_8_0_t121[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t123 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_8_0_t124 = FSM_dct_8x8_stage_8_0_t123[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t125 = FSM_dct_8x8_stage_8_0_t124[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t126 = i_data_in[FSM_dct_8x8_stage_8_0_t125 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t127 = FSM_dct_8x8_stage_8_0_t119;
    FSM_dct_8x8_stage_8_0_t127[FSM_dct_8x8_stage_8_0_t122 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t126;
    FSM_dct_8x8_stage_8_0_t128 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_8_0_t129 = FSM_dct_8x8_stage_8_0_t128[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t130 = FSM_dct_8x8_stage_8_0_t129[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t131 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_8_0_t132 = FSM_dct_8x8_stage_8_0_t131[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t133 = FSM_dct_8x8_stage_8_0_t132[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t134 = i_data_in[FSM_dct_8x8_stage_8_0_t133 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t135 = FSM_dct_8x8_stage_8_0_t127;
    FSM_dct_8x8_stage_8_0_t135[FSM_dct_8x8_stage_8_0_t130 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t134;
    FSM_dct_8x8_stage_8_0_t136 = 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_8_0_t137 = FSM_dct_8x8_stage_8_0_t136[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t138 = 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_8_0_t139 = FSM_dct_8x8_stage_8_0_t138[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t140 = i_data_in[FSM_dct_8x8_stage_8_0_t139 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t141 = FSM_dct_8x8_stage_8_0_t135;
    FSM_dct_8x8_stage_8_0_t141[FSM_dct_8x8_stage_8_0_t137 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t140;
    FSM_dct_8x8_stage_8_0_t142 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_8_0_t143 = FSM_dct_8x8_stage_8_0_t142[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t144 = FSM_dct_8x8_stage_8_0_t143[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t145 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_8_0_t146 = FSM_dct_8x8_stage_8_0_t145[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t147 = FSM_dct_8x8_stage_8_0_t146[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t148 = i_data_in[FSM_dct_8x8_stage_8_0_t147 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t149 = FSM_dct_8x8_stage_8_0_t141;
    FSM_dct_8x8_stage_8_0_t149[FSM_dct_8x8_stage_8_0_t144 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t148;
    FSM_dct_8x8_stage_8_0_t150 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_8_0_t151 = FSM_dct_8x8_stage_8_0_t150[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t152 = FSM_dct_8x8_stage_8_0_t151[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t153 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_8_0_t154 = FSM_dct_8x8_stage_8_0_t153[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t155 = FSM_dct_8x8_stage_8_0_t154[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t156 = i_data_in[FSM_dct_8x8_stage_8_0_t155 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t157 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_8_0_t158 = FSM_dct_8x8_stage_8_0_t157[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t159 = FSM_dct_8x8_stage_8_0_t158[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t160 = i_data_in[FSM_dct_8x8_stage_8_0_t159 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t161 = FSM_dct_8x8_stage_8_0_t156 + FSM_dct_8x8_stage_8_0_t160;
    FSM_dct_8x8_stage_8_0_t162 = FSM_dct_8x8_stage_8_0_t161[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t163 = FSM_dct_8x8_stage_8_0_t149;
    FSM_dct_8x8_stage_8_0_t163[FSM_dct_8x8_stage_8_0_t152 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t162;
    FSM_dct_8x8_stage_8_0_t164 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_8_0_t165 = FSM_dct_8x8_stage_8_0_t164[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t166 = FSM_dct_8x8_stage_8_0_t165[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t167 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_8_0_t168 = FSM_dct_8x8_stage_8_0_t167[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t169 = FSM_dct_8x8_stage_8_0_t168[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t170 = i_data_in[FSM_dct_8x8_stage_8_0_t169 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t171 = FSM_dct_8x8_stage_8_0_t163;
    FSM_dct_8x8_stage_8_0_t171[FSM_dct_8x8_stage_8_0_t166 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t170;
    FSM_dct_8x8_stage_8_0_t172 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_8_0_t173 = FSM_dct_8x8_stage_8_0_t172[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t174 = FSM_dct_8x8_stage_8_0_t173[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t175 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_8_0_t176 = FSM_dct_8x8_stage_8_0_t175[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t177 = FSM_dct_8x8_stage_8_0_t176[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t178 = i_data_in[FSM_dct_8x8_stage_8_0_t177 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t179 = FSM_dct_8x8_stage_8_0_t171;
    FSM_dct_8x8_stage_8_0_t179[FSM_dct_8x8_stage_8_0_t174 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t178;
    FSM_dct_8x8_stage_8_0_t180 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_8_0_t181 = FSM_dct_8x8_stage_8_0_t180[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t182 = FSM_dct_8x8_stage_8_0_t181[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t183 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_8_0_t184 = FSM_dct_8x8_stage_8_0_t183[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t185 = FSM_dct_8x8_stage_8_0_t184[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t186 = i_data_in[FSM_dct_8x8_stage_8_0_t185 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t187 = FSM_dct_8x8_stage_8_0_t179;
    FSM_dct_8x8_stage_8_0_t187[FSM_dct_8x8_stage_8_0_t182 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t186;
    FSM_dct_8x8_stage_8_0_t188 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_8_0_t189 = FSM_dct_8x8_stage_8_0_t188[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t190 = FSM_dct_8x8_stage_8_0_t189[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t191 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_8_0_t192 = FSM_dct_8x8_stage_8_0_t191[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t193 = FSM_dct_8x8_stage_8_0_t192[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t194 = i_data_in[FSM_dct_8x8_stage_8_0_t193 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t195 = FSM_dct_8x8_stage_8_0_t187;
    FSM_dct_8x8_stage_8_0_t195[FSM_dct_8x8_stage_8_0_t190 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t194;
    FSM_dct_8x8_stage_8_0_t196 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_8_0_t197 = FSM_dct_8x8_stage_8_0_t196[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t198 = FSM_dct_8x8_stage_8_0_t197[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t199 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_8_0_t200 = FSM_dct_8x8_stage_8_0_t199[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t201 = FSM_dct_8x8_stage_8_0_t200[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t202 = i_data_in[FSM_dct_8x8_stage_8_0_t201 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t203 = FSM_dct_8x8_stage_8_0_t195;
    FSM_dct_8x8_stage_8_0_t203[FSM_dct_8x8_stage_8_0_t198 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t202;
    FSM_dct_8x8_stage_8_0_t204 = 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_8_0_t205 = FSM_dct_8x8_stage_8_0_t204[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t206 = 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_8_0_t207 = FSM_dct_8x8_stage_8_0_t206[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t208 = i_data_in[FSM_dct_8x8_stage_8_0_t207 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t209 = FSM_dct_8x8_stage_8_0_t203;
    FSM_dct_8x8_stage_8_0_t209[FSM_dct_8x8_stage_8_0_t205 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t208;
    FSM_dct_8x8_stage_8_0_t210 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_8_0_t211 = FSM_dct_8x8_stage_8_0_t210[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t212 = FSM_dct_8x8_stage_8_0_t211[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t213 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_8_0_t214 = FSM_dct_8x8_stage_8_0_t213[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t215 = FSM_dct_8x8_stage_8_0_t214[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t216 = i_data_in[FSM_dct_8x8_stage_8_0_t215 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t217 = FSM_dct_8x8_stage_8_0_t209;
    FSM_dct_8x8_stage_8_0_t217[FSM_dct_8x8_stage_8_0_t212 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t216;
    FSM_dct_8x8_stage_8_0_t218 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_8_0_t219 = FSM_dct_8x8_stage_8_0_t218[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t220 = FSM_dct_8x8_stage_8_0_t219[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t221 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_8_0_t222 = FSM_dct_8x8_stage_8_0_t221[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t223 = FSM_dct_8x8_stage_8_0_t222[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t224 = i_data_in[FSM_dct_8x8_stage_8_0_t223 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t225 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_8_0_t226 = FSM_dct_8x8_stage_8_0_t225[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t227 = FSM_dct_8x8_stage_8_0_t226[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t228 = i_data_in[FSM_dct_8x8_stage_8_0_t227 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t229 = FSM_dct_8x8_stage_8_0_t224 + FSM_dct_8x8_stage_8_0_t228;
    FSM_dct_8x8_stage_8_0_t230 = FSM_dct_8x8_stage_8_0_t229[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t231 = FSM_dct_8x8_stage_8_0_t217;
    FSM_dct_8x8_stage_8_0_t231[FSM_dct_8x8_stage_8_0_t220 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t230;
    FSM_dct_8x8_stage_8_0_t232 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_8_0_t233 = FSM_dct_8x8_stage_8_0_t232[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t234 = FSM_dct_8x8_stage_8_0_t233[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t235 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_8_0_t236 = FSM_dct_8x8_stage_8_0_t235[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t237 = FSM_dct_8x8_stage_8_0_t236[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t238 = i_data_in[FSM_dct_8x8_stage_8_0_t237 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t239 = FSM_dct_8x8_stage_8_0_t231;
    FSM_dct_8x8_stage_8_0_t239[FSM_dct_8x8_stage_8_0_t234 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t238;
    FSM_dct_8x8_stage_8_0_t240 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_8_0_t241 = FSM_dct_8x8_stage_8_0_t240[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t242 = FSM_dct_8x8_stage_8_0_t241[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t243 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_8_0_t244 = FSM_dct_8x8_stage_8_0_t243[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t245 = FSM_dct_8x8_stage_8_0_t244[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t246 = i_data_in[FSM_dct_8x8_stage_8_0_t245 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t247 = FSM_dct_8x8_stage_8_0_t239;
    FSM_dct_8x8_stage_8_0_t247[FSM_dct_8x8_stage_8_0_t242 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t246;
    FSM_dct_8x8_stage_8_0_t248 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_8_0_t249 = FSM_dct_8x8_stage_8_0_t248[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t250 = FSM_dct_8x8_stage_8_0_t249[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t251 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_8_0_t252 = FSM_dct_8x8_stage_8_0_t251[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t253 = FSM_dct_8x8_stage_8_0_t252[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t254 = i_data_in[FSM_dct_8x8_stage_8_0_t253 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t255 = FSM_dct_8x8_stage_8_0_t247;
    FSM_dct_8x8_stage_8_0_t255[FSM_dct_8x8_stage_8_0_t250 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t254;
    FSM_dct_8x8_stage_8_0_t256 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_8_0_t257 = FSM_dct_8x8_stage_8_0_t256[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t258 = FSM_dct_8x8_stage_8_0_t257[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t259 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_8_0_t260 = FSM_dct_8x8_stage_8_0_t259[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t261 = FSM_dct_8x8_stage_8_0_t260[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t262 = i_data_in[FSM_dct_8x8_stage_8_0_t261 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t263 = FSM_dct_8x8_stage_8_0_t255;
    FSM_dct_8x8_stage_8_0_t263[FSM_dct_8x8_stage_8_0_t258 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t262;
    FSM_dct_8x8_stage_8_0_t264 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_8_0_t265 = FSM_dct_8x8_stage_8_0_t264[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t266 = FSM_dct_8x8_stage_8_0_t265[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t267 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_8_0_t268 = FSM_dct_8x8_stage_8_0_t267[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t269 = FSM_dct_8x8_stage_8_0_t268[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t270 = i_data_in[FSM_dct_8x8_stage_8_0_t269 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t271 = FSM_dct_8x8_stage_8_0_t263;
    FSM_dct_8x8_stage_8_0_t271[FSM_dct_8x8_stage_8_0_t266 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t270;
    FSM_dct_8x8_stage_8_0_t272 = 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_8_0_t273 = FSM_dct_8x8_stage_8_0_t272[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t274 = 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_8_0_t275 = FSM_dct_8x8_stage_8_0_t274[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t276 = i_data_in[FSM_dct_8x8_stage_8_0_t275 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t277 = FSM_dct_8x8_stage_8_0_t271;
    FSM_dct_8x8_stage_8_0_t277[FSM_dct_8x8_stage_8_0_t273 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t276;
    FSM_dct_8x8_stage_8_0_t278 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_8_0_t279 = FSM_dct_8x8_stage_8_0_t278[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t280 = FSM_dct_8x8_stage_8_0_t279[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t281 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_8_0_t282 = FSM_dct_8x8_stage_8_0_t281[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t283 = FSM_dct_8x8_stage_8_0_t282[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t284 = i_data_in[FSM_dct_8x8_stage_8_0_t283 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t285 = FSM_dct_8x8_stage_8_0_t277;
    FSM_dct_8x8_stage_8_0_t285[FSM_dct_8x8_stage_8_0_t280 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t284;
    FSM_dct_8x8_stage_8_0_t286 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_8_0_t287 = FSM_dct_8x8_stage_8_0_t286[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t288 = FSM_dct_8x8_stage_8_0_t287[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t289 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_8_0_t290 = FSM_dct_8x8_stage_8_0_t289[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t291 = FSM_dct_8x8_stage_8_0_t290[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t292 = i_data_in[FSM_dct_8x8_stage_8_0_t291 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t293 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_8_0_t294 = FSM_dct_8x8_stage_8_0_t293[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t295 = FSM_dct_8x8_stage_8_0_t294[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t296 = i_data_in[FSM_dct_8x8_stage_8_0_t295 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t297 = FSM_dct_8x8_stage_8_0_t292 + FSM_dct_8x8_stage_8_0_t296;
    FSM_dct_8x8_stage_8_0_t298 = FSM_dct_8x8_stage_8_0_t297[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t299 = FSM_dct_8x8_stage_8_0_t285;
    FSM_dct_8x8_stage_8_0_t299[FSM_dct_8x8_stage_8_0_t288 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t298;
    FSM_dct_8x8_stage_8_0_t300 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_8_0_t301 = FSM_dct_8x8_stage_8_0_t300[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t302 = FSM_dct_8x8_stage_8_0_t301[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t303 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_8_0_t304 = FSM_dct_8x8_stage_8_0_t303[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t305 = FSM_dct_8x8_stage_8_0_t304[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t306 = i_data_in[FSM_dct_8x8_stage_8_0_t305 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t307 = FSM_dct_8x8_stage_8_0_t299;
    FSM_dct_8x8_stage_8_0_t307[FSM_dct_8x8_stage_8_0_t302 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t306;
    FSM_dct_8x8_stage_8_0_t308 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_8_0_t309 = FSM_dct_8x8_stage_8_0_t308[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t310 = FSM_dct_8x8_stage_8_0_t309[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t311 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_8_0_t312 = FSM_dct_8x8_stage_8_0_t311[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t313 = FSM_dct_8x8_stage_8_0_t312[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t314 = i_data_in[FSM_dct_8x8_stage_8_0_t313 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t315 = FSM_dct_8x8_stage_8_0_t307;
    FSM_dct_8x8_stage_8_0_t315[FSM_dct_8x8_stage_8_0_t310 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t314;
    FSM_dct_8x8_stage_8_0_t316 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_8_0_t317 = FSM_dct_8x8_stage_8_0_t316[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t318 = FSM_dct_8x8_stage_8_0_t317[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t319 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_8_0_t320 = FSM_dct_8x8_stage_8_0_t319[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t321 = FSM_dct_8x8_stage_8_0_t320[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t322 = i_data_in[FSM_dct_8x8_stage_8_0_t321 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t323 = FSM_dct_8x8_stage_8_0_t315;
    FSM_dct_8x8_stage_8_0_t323[FSM_dct_8x8_stage_8_0_t318 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t322;
    FSM_dct_8x8_stage_8_0_t324 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_8_0_t325 = FSM_dct_8x8_stage_8_0_t324[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t326 = FSM_dct_8x8_stage_8_0_t325[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t327 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_8_0_t328 = FSM_dct_8x8_stage_8_0_t327[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t329 = FSM_dct_8x8_stage_8_0_t328[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t330 = i_data_in[FSM_dct_8x8_stage_8_0_t329 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t331 = FSM_dct_8x8_stage_8_0_t323;
    FSM_dct_8x8_stage_8_0_t331[FSM_dct_8x8_stage_8_0_t326 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t330;
    FSM_dct_8x8_stage_8_0_t332 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_8_0_t333 = FSM_dct_8x8_stage_8_0_t332[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t334 = FSM_dct_8x8_stage_8_0_t333[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t335 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_8_0_t336 = FSM_dct_8x8_stage_8_0_t335[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t337 = FSM_dct_8x8_stage_8_0_t336[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t338 = i_data_in[FSM_dct_8x8_stage_8_0_t337 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t339 = FSM_dct_8x8_stage_8_0_t331;
    FSM_dct_8x8_stage_8_0_t339[FSM_dct_8x8_stage_8_0_t334 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t338;
    FSM_dct_8x8_stage_8_0_t340 = 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_8_0_t341 = FSM_dct_8x8_stage_8_0_t340[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t342 = 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_8_0_t343 = FSM_dct_8x8_stage_8_0_t342[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t344 = i_data_in[FSM_dct_8x8_stage_8_0_t343 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t345 = FSM_dct_8x8_stage_8_0_t339;
    FSM_dct_8x8_stage_8_0_t345[FSM_dct_8x8_stage_8_0_t341 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t344;
    FSM_dct_8x8_stage_8_0_t346 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_8_0_t347 = FSM_dct_8x8_stage_8_0_t346[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t348 = FSM_dct_8x8_stage_8_0_t347[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t349 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_8_0_t350 = FSM_dct_8x8_stage_8_0_t349[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t351 = FSM_dct_8x8_stage_8_0_t350[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t352 = i_data_in[FSM_dct_8x8_stage_8_0_t351 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t353 = FSM_dct_8x8_stage_8_0_t345;
    FSM_dct_8x8_stage_8_0_t353[FSM_dct_8x8_stage_8_0_t348 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t352;
    FSM_dct_8x8_stage_8_0_t354 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_8_0_t355 = FSM_dct_8x8_stage_8_0_t354[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t356 = FSM_dct_8x8_stage_8_0_t355[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t357 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_8_0_t358 = FSM_dct_8x8_stage_8_0_t357[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t359 = FSM_dct_8x8_stage_8_0_t358[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t360 = i_data_in[FSM_dct_8x8_stage_8_0_t359 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t361 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_8_0_t362 = FSM_dct_8x8_stage_8_0_t361[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t363 = FSM_dct_8x8_stage_8_0_t362[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t364 = i_data_in[FSM_dct_8x8_stage_8_0_t363 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t365 = FSM_dct_8x8_stage_8_0_t360 + FSM_dct_8x8_stage_8_0_t364;
    FSM_dct_8x8_stage_8_0_t366 = FSM_dct_8x8_stage_8_0_t365[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t367 = FSM_dct_8x8_stage_8_0_t353;
    FSM_dct_8x8_stage_8_0_t367[FSM_dct_8x8_stage_8_0_t356 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t366;
    FSM_dct_8x8_stage_8_0_t368 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_8_0_t369 = FSM_dct_8x8_stage_8_0_t368[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t370 = FSM_dct_8x8_stage_8_0_t369[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t371 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_8_0_t372 = FSM_dct_8x8_stage_8_0_t371[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t373 = FSM_dct_8x8_stage_8_0_t372[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t374 = i_data_in[FSM_dct_8x8_stage_8_0_t373 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t375 = FSM_dct_8x8_stage_8_0_t367;
    FSM_dct_8x8_stage_8_0_t375[FSM_dct_8x8_stage_8_0_t370 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t374;
    FSM_dct_8x8_stage_8_0_t376 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_8_0_t377 = FSM_dct_8x8_stage_8_0_t376[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t378 = FSM_dct_8x8_stage_8_0_t377[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t379 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_8_0_t380 = FSM_dct_8x8_stage_8_0_t379[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t381 = FSM_dct_8x8_stage_8_0_t380[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t382 = i_data_in[FSM_dct_8x8_stage_8_0_t381 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t383 = FSM_dct_8x8_stage_8_0_t375;
    FSM_dct_8x8_stage_8_0_t383[FSM_dct_8x8_stage_8_0_t378 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t382;
    FSM_dct_8x8_stage_8_0_t384 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_8_0_t385 = FSM_dct_8x8_stage_8_0_t384[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t386 = FSM_dct_8x8_stage_8_0_t385[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t387 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_8_0_t388 = FSM_dct_8x8_stage_8_0_t387[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t389 = FSM_dct_8x8_stage_8_0_t388[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t390 = i_data_in[FSM_dct_8x8_stage_8_0_t389 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t391 = FSM_dct_8x8_stage_8_0_t383;
    FSM_dct_8x8_stage_8_0_t391[FSM_dct_8x8_stage_8_0_t386 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t390;
    FSM_dct_8x8_stage_8_0_t392 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_8_0_t393 = FSM_dct_8x8_stage_8_0_t392[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t394 = FSM_dct_8x8_stage_8_0_t393[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t395 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_8_0_t396 = FSM_dct_8x8_stage_8_0_t395[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t397 = FSM_dct_8x8_stage_8_0_t396[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t398 = i_data_in[FSM_dct_8x8_stage_8_0_t397 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t399 = FSM_dct_8x8_stage_8_0_t391;
    FSM_dct_8x8_stage_8_0_t399[FSM_dct_8x8_stage_8_0_t394 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t398;
    FSM_dct_8x8_stage_8_0_t400 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_8_0_t401 = FSM_dct_8x8_stage_8_0_t400[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t402 = FSM_dct_8x8_stage_8_0_t401[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t403 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_8_0_t404 = FSM_dct_8x8_stage_8_0_t403[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t405 = FSM_dct_8x8_stage_8_0_t404[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t406 = i_data_in[FSM_dct_8x8_stage_8_0_t405 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t407 = FSM_dct_8x8_stage_8_0_t399;
    FSM_dct_8x8_stage_8_0_t407[FSM_dct_8x8_stage_8_0_t402 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t406;
    FSM_dct_8x8_stage_8_0_t408 = 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_8_0_t409 = FSM_dct_8x8_stage_8_0_t408[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t410 = 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_8_0_t411 = FSM_dct_8x8_stage_8_0_t410[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t412 = i_data_in[FSM_dct_8x8_stage_8_0_t411 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t413 = FSM_dct_8x8_stage_8_0_t407;
    FSM_dct_8x8_stage_8_0_t413[FSM_dct_8x8_stage_8_0_t409 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t412;
    FSM_dct_8x8_stage_8_0_t414 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_8_0_t415 = FSM_dct_8x8_stage_8_0_t414[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t416 = FSM_dct_8x8_stage_8_0_t415[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t417 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_8_0_t418 = FSM_dct_8x8_stage_8_0_t417[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t419 = FSM_dct_8x8_stage_8_0_t418[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t420 = i_data_in[FSM_dct_8x8_stage_8_0_t419 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t421 = FSM_dct_8x8_stage_8_0_t413;
    FSM_dct_8x8_stage_8_0_t421[FSM_dct_8x8_stage_8_0_t416 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t420;
    FSM_dct_8x8_stage_8_0_t422 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_8_0_t423 = FSM_dct_8x8_stage_8_0_t422[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t424 = FSM_dct_8x8_stage_8_0_t423[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t425 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_8_0_t426 = FSM_dct_8x8_stage_8_0_t425[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t427 = FSM_dct_8x8_stage_8_0_t426[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t428 = i_data_in[FSM_dct_8x8_stage_8_0_t427 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t429 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_8_0_t430 = FSM_dct_8x8_stage_8_0_t429[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t431 = FSM_dct_8x8_stage_8_0_t430[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t432 = i_data_in[FSM_dct_8x8_stage_8_0_t431 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t433 = FSM_dct_8x8_stage_8_0_t428 + FSM_dct_8x8_stage_8_0_t432;
    FSM_dct_8x8_stage_8_0_t434 = FSM_dct_8x8_stage_8_0_t433[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t435 = FSM_dct_8x8_stage_8_0_t421;
    FSM_dct_8x8_stage_8_0_t435[FSM_dct_8x8_stage_8_0_t424 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t434;
    FSM_dct_8x8_stage_8_0_t436 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_8_0_t437 = FSM_dct_8x8_stage_8_0_t436[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t438 = FSM_dct_8x8_stage_8_0_t437[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t439 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_8_0_t440 = FSM_dct_8x8_stage_8_0_t439[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t441 = FSM_dct_8x8_stage_8_0_t440[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t442 = i_data_in[FSM_dct_8x8_stage_8_0_t441 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t443 = FSM_dct_8x8_stage_8_0_t435;
    FSM_dct_8x8_stage_8_0_t443[FSM_dct_8x8_stage_8_0_t438 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t442;
    FSM_dct_8x8_stage_8_0_t444 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_8_0_t445 = FSM_dct_8x8_stage_8_0_t444[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t446 = FSM_dct_8x8_stage_8_0_t445[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t447 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_8_0_t448 = FSM_dct_8x8_stage_8_0_t447[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t449 = FSM_dct_8x8_stage_8_0_t448[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t450 = i_data_in[FSM_dct_8x8_stage_8_0_t449 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t451 = FSM_dct_8x8_stage_8_0_t443;
    FSM_dct_8x8_stage_8_0_t451[FSM_dct_8x8_stage_8_0_t446 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t450;
    FSM_dct_8x8_stage_8_0_t452 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_8_0_t453 = FSM_dct_8x8_stage_8_0_t452[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t454 = FSM_dct_8x8_stage_8_0_t453[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t455 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_8_0_t456 = FSM_dct_8x8_stage_8_0_t455[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t457 = FSM_dct_8x8_stage_8_0_t456[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t458 = i_data_in[FSM_dct_8x8_stage_8_0_t457 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t459 = FSM_dct_8x8_stage_8_0_t451;
    FSM_dct_8x8_stage_8_0_t459[FSM_dct_8x8_stage_8_0_t454 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t458;
    FSM_dct_8x8_stage_8_0_t460 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_8_0_t461 = FSM_dct_8x8_stage_8_0_t460[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t462 = FSM_dct_8x8_stage_8_0_t461[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t463 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_8_0_t464 = FSM_dct_8x8_stage_8_0_t463[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t465 = FSM_dct_8x8_stage_8_0_t464[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t466 = i_data_in[FSM_dct_8x8_stage_8_0_t465 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t467 = FSM_dct_8x8_stage_8_0_t459;
    FSM_dct_8x8_stage_8_0_t467[FSM_dct_8x8_stage_8_0_t462 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t466;
    FSM_dct_8x8_stage_8_0_t468 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_8_0_t469 = FSM_dct_8x8_stage_8_0_t468[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t470 = FSM_dct_8x8_stage_8_0_t469[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t471 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_8_0_t472 = FSM_dct_8x8_stage_8_0_t471[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t473 = FSM_dct_8x8_stage_8_0_t472[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t474 = i_data_in[FSM_dct_8x8_stage_8_0_t473 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t475 = FSM_dct_8x8_stage_8_0_t467;
    FSM_dct_8x8_stage_8_0_t475[FSM_dct_8x8_stage_8_0_t470 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t474;
    FSM_dct_8x8_stage_8_0_t476 = 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_8_0_t477 = FSM_dct_8x8_stage_8_0_t476[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t478 = 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_8_0_t479 = FSM_dct_8x8_stage_8_0_t478[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t480 = i_data_in[FSM_dct_8x8_stage_8_0_t479 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t481 = FSM_dct_8x8_stage_8_0_t475;
    FSM_dct_8x8_stage_8_0_t481[FSM_dct_8x8_stage_8_0_t477 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t480;
    FSM_dct_8x8_stage_8_0_t482 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_8_0_t483 = FSM_dct_8x8_stage_8_0_t482[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t484 = FSM_dct_8x8_stage_8_0_t483[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t485 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_8_0_t486 = FSM_dct_8x8_stage_8_0_t485[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t487 = FSM_dct_8x8_stage_8_0_t486[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t488 = i_data_in[FSM_dct_8x8_stage_8_0_t487 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t489 = FSM_dct_8x8_stage_8_0_t481;
    FSM_dct_8x8_stage_8_0_t489[FSM_dct_8x8_stage_8_0_t484 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t488;
    FSM_dct_8x8_stage_8_0_t490 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_8_0_t491 = FSM_dct_8x8_stage_8_0_t490[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t492 = FSM_dct_8x8_stage_8_0_t491[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t493 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_8_0_t494 = FSM_dct_8x8_stage_8_0_t493[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t495 = FSM_dct_8x8_stage_8_0_t494[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t496 = i_data_in[FSM_dct_8x8_stage_8_0_t495 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t497 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_8_0_t498 = FSM_dct_8x8_stage_8_0_t497[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t499 = FSM_dct_8x8_stage_8_0_t498[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t500 = i_data_in[FSM_dct_8x8_stage_8_0_t499 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t501 = FSM_dct_8x8_stage_8_0_t496 + FSM_dct_8x8_stage_8_0_t500;
    FSM_dct_8x8_stage_8_0_t502 = FSM_dct_8x8_stage_8_0_t501[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t503 = FSM_dct_8x8_stage_8_0_t489;
    FSM_dct_8x8_stage_8_0_t503[FSM_dct_8x8_stage_8_0_t492 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t502;
    FSM_dct_8x8_stage_8_0_t504 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_8_0_t505 = FSM_dct_8x8_stage_8_0_t504[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t506 = FSM_dct_8x8_stage_8_0_t505[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t507 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_8_0_t508 = FSM_dct_8x8_stage_8_0_t507[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t509 = FSM_dct_8x8_stage_8_0_t508[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t510 = i_data_in[FSM_dct_8x8_stage_8_0_t509 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t511 = FSM_dct_8x8_stage_8_0_t503;
    FSM_dct_8x8_stage_8_0_t511[FSM_dct_8x8_stage_8_0_t506 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t510;
    FSM_dct_8x8_stage_8_0_t512 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_8_0_t513 = FSM_dct_8x8_stage_8_0_t512[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t514 = FSM_dct_8x8_stage_8_0_t513[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t515 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_8_0_t516 = FSM_dct_8x8_stage_8_0_t515[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t517 = FSM_dct_8x8_stage_8_0_t516[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t518 = i_data_in[FSM_dct_8x8_stage_8_0_t517 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t519 = FSM_dct_8x8_stage_8_0_t511;
    FSM_dct_8x8_stage_8_0_t519[FSM_dct_8x8_stage_8_0_t514 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t518;
    FSM_dct_8x8_stage_8_0_t520 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_8_0_t521 = FSM_dct_8x8_stage_8_0_t520[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t522 = FSM_dct_8x8_stage_8_0_t521[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t523 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_8_0_t524 = FSM_dct_8x8_stage_8_0_t523[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t525 = FSM_dct_8x8_stage_8_0_t524[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t526 = i_data_in[FSM_dct_8x8_stage_8_0_t525 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t527 = FSM_dct_8x8_stage_8_0_t519;
    FSM_dct_8x8_stage_8_0_t527[FSM_dct_8x8_stage_8_0_t522 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t526;
    FSM_dct_8x8_stage_8_0_t528 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_8_0_t529 = FSM_dct_8x8_stage_8_0_t528[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t530 = FSM_dct_8x8_stage_8_0_t529[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t531 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_8_0_t532 = FSM_dct_8x8_stage_8_0_t531[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t533 = FSM_dct_8x8_stage_8_0_t532[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t534 = i_data_in[FSM_dct_8x8_stage_8_0_t533 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t535 = FSM_dct_8x8_stage_8_0_t527;
    FSM_dct_8x8_stage_8_0_t535[FSM_dct_8x8_stage_8_0_t530 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t534;
    FSM_dct_8x8_stage_8_0_t536 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_8_0_t537 = FSM_dct_8x8_stage_8_0_t536[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t538 = FSM_dct_8x8_stage_8_0_t537[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t539 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_8_0_t540 = FSM_dct_8x8_stage_8_0_t539[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t541 = FSM_dct_8x8_stage_8_0_t540[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t542 = i_data_in[FSM_dct_8x8_stage_8_0_t541 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t543 = FSM_dct_8x8_stage_8_0_t535;
    FSM_dct_8x8_stage_8_0_t543[FSM_dct_8x8_stage_8_0_t538 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t542;
end

always @* begin
    FSM_dct_8x8_stage_8_0_t0 = 32'b0;
    FSM_dct_8x8_stage_8_0_t1 = FSM_dct_8x8_stage_8_0_t0[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t2 = 32'b0;
    FSM_dct_8x8_stage_8_0_t3 = FSM_dct_8x8_stage_8_0_t2[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t4 = i_data_in[FSM_dct_8x8_stage_8_0_t3 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t5 = 2048'b0;
    FSM_dct_8x8_stage_8_0_t5[FSM_dct_8x8_stage_8_0_t1 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t4;
    FSM_dct_8x8_stage_8_0_t6 = 32'b00000000000000000000000000001000 + 32'b0;
    FSM_dct_8x8_stage_8_0_t7 = FSM_dct_8x8_stage_8_0_t6[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t8 = FSM_dct_8x8_stage_8_0_t7[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t9 = 32'b00000000000000000000000000001000 + 32'b0;
    FSM_dct_8x8_stage_8_0_t10 = FSM_dct_8x8_stage_8_0_t9[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t11 = FSM_dct_8x8_stage_8_0_t10[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t12 = i_data_in[FSM_dct_8x8_stage_8_0_t11 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t13 = FSM_dct_8x8_stage_8_0_t5;
    FSM_dct_8x8_stage_8_0_t13[FSM_dct_8x8_stage_8_0_t8 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t12;
    FSM_dct_8x8_stage_8_0_t14 = 32'b00000000000000000000000000010000 + 32'b0;
    FSM_dct_8x8_stage_8_0_t15 = FSM_dct_8x8_stage_8_0_t14[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t16 = FSM_dct_8x8_stage_8_0_t15[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t17 = 32'b00000000000000000000000000010000 + 32'b0;
    FSM_dct_8x8_stage_8_0_t18 = FSM_dct_8x8_stage_8_0_t17[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t19 = FSM_dct_8x8_stage_8_0_t18[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t20 = i_data_in[FSM_dct_8x8_stage_8_0_t19 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t21 = 32'b00000000000000000000000000011000 + 32'b0;
    FSM_dct_8x8_stage_8_0_t22 = FSM_dct_8x8_stage_8_0_t21[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t23 = FSM_dct_8x8_stage_8_0_t22[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t24 = i_data_in[FSM_dct_8x8_stage_8_0_t23 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t25 = FSM_dct_8x8_stage_8_0_t20 + FSM_dct_8x8_stage_8_0_t24;
    FSM_dct_8x8_stage_8_0_t26 = FSM_dct_8x8_stage_8_0_t25[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t27 = FSM_dct_8x8_stage_8_0_t13;
    FSM_dct_8x8_stage_8_0_t27[FSM_dct_8x8_stage_8_0_t16 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t26;
    FSM_dct_8x8_stage_8_0_t28 = 32'b00000000000000000000000000011000 + 32'b0;
    FSM_dct_8x8_stage_8_0_t29 = FSM_dct_8x8_stage_8_0_t28[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t30 = FSM_dct_8x8_stage_8_0_t29[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t31 = 32'b00000000000000000000000000011000 + 32'b0;
    FSM_dct_8x8_stage_8_0_t32 = FSM_dct_8x8_stage_8_0_t31[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t33 = FSM_dct_8x8_stage_8_0_t32[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t34 = i_data_in[FSM_dct_8x8_stage_8_0_t33 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t35 = FSM_dct_8x8_stage_8_0_t27;
    FSM_dct_8x8_stage_8_0_t35[FSM_dct_8x8_stage_8_0_t30 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t34;
    FSM_dct_8x8_stage_8_0_t36 = 32'b00000000000000000000000000100000 + 32'b0;
    FSM_dct_8x8_stage_8_0_t37 = FSM_dct_8x8_stage_8_0_t36[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t38 = FSM_dct_8x8_stage_8_0_t37[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t39 = 32'b00000000000000000000000000100000 + 32'b0;
    FSM_dct_8x8_stage_8_0_t40 = FSM_dct_8x8_stage_8_0_t39[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t41 = FSM_dct_8x8_stage_8_0_t40[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t42 = i_data_in[FSM_dct_8x8_stage_8_0_t41 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t43 = FSM_dct_8x8_stage_8_0_t35;
    FSM_dct_8x8_stage_8_0_t43[FSM_dct_8x8_stage_8_0_t38 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t42;
    FSM_dct_8x8_stage_8_0_t44 = 32'b00000000000000000000000000101000 + 32'b0;
    FSM_dct_8x8_stage_8_0_t45 = FSM_dct_8x8_stage_8_0_t44[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t46 = FSM_dct_8x8_stage_8_0_t45[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t47 = 32'b00000000000000000000000000101000 + 32'b0;
    FSM_dct_8x8_stage_8_0_t48 = FSM_dct_8x8_stage_8_0_t47[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t49 = FSM_dct_8x8_stage_8_0_t48[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t50 = i_data_in[FSM_dct_8x8_stage_8_0_t49 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t51 = FSM_dct_8x8_stage_8_0_t43;
    FSM_dct_8x8_stage_8_0_t51[FSM_dct_8x8_stage_8_0_t46 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t50;
    FSM_dct_8x8_stage_8_0_t52 = 32'b00000000000000000000000000110000 + 32'b0;
    FSM_dct_8x8_stage_8_0_t53 = FSM_dct_8x8_stage_8_0_t52[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t54 = FSM_dct_8x8_stage_8_0_t53[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t55 = 32'b00000000000000000000000000110000 + 32'b0;
    FSM_dct_8x8_stage_8_0_t56 = FSM_dct_8x8_stage_8_0_t55[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t57 = FSM_dct_8x8_stage_8_0_t56[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t58 = i_data_in[FSM_dct_8x8_stage_8_0_t57 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t59 = FSM_dct_8x8_stage_8_0_t51;
    FSM_dct_8x8_stage_8_0_t59[FSM_dct_8x8_stage_8_0_t54 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t58;
    FSM_dct_8x8_stage_8_0_t60 = 32'b00000000000000000000000000111000 + 32'b0;
    FSM_dct_8x8_stage_8_0_t61 = FSM_dct_8x8_stage_8_0_t60[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t62 = FSM_dct_8x8_stage_8_0_t61[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t63 = 32'b00000000000000000000000000111000 + 32'b0;
    FSM_dct_8x8_stage_8_0_t64 = FSM_dct_8x8_stage_8_0_t63[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t65 = FSM_dct_8x8_stage_8_0_t64[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t66 = i_data_in[FSM_dct_8x8_stage_8_0_t65 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t67 = FSM_dct_8x8_stage_8_0_t59;
    FSM_dct_8x8_stage_8_0_t67[FSM_dct_8x8_stage_8_0_t62 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t66;
    FSM_dct_8x8_stage_8_0_t68 = 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_8_0_t69 = FSM_dct_8x8_stage_8_0_t68[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t70 = 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_8_0_t71 = FSM_dct_8x8_stage_8_0_t70[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t72 = i_data_in[FSM_dct_8x8_stage_8_0_t71 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t73 = FSM_dct_8x8_stage_8_0_t67;
    FSM_dct_8x8_stage_8_0_t73[FSM_dct_8x8_stage_8_0_t69 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t72;
    FSM_dct_8x8_stage_8_0_t74 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_8_0_t75 = FSM_dct_8x8_stage_8_0_t74[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t76 = FSM_dct_8x8_stage_8_0_t75[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t77 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_8_0_t78 = FSM_dct_8x8_stage_8_0_t77[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t79 = FSM_dct_8x8_stage_8_0_t78[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t80 = i_data_in[FSM_dct_8x8_stage_8_0_t79 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t81 = FSM_dct_8x8_stage_8_0_t73;
    FSM_dct_8x8_stage_8_0_t81[FSM_dct_8x8_stage_8_0_t76 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t80;
    FSM_dct_8x8_stage_8_0_t82 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_8_0_t83 = FSM_dct_8x8_stage_8_0_t82[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t84 = FSM_dct_8x8_stage_8_0_t83[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t85 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_8_0_t86 = FSM_dct_8x8_stage_8_0_t85[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t87 = FSM_dct_8x8_stage_8_0_t86[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t88 = i_data_in[FSM_dct_8x8_stage_8_0_t87 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t89 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_8_0_t90 = FSM_dct_8x8_stage_8_0_t89[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t91 = FSM_dct_8x8_stage_8_0_t90[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t92 = i_data_in[FSM_dct_8x8_stage_8_0_t91 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t93 = FSM_dct_8x8_stage_8_0_t88 + FSM_dct_8x8_stage_8_0_t92;
    FSM_dct_8x8_stage_8_0_t94 = FSM_dct_8x8_stage_8_0_t93[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t95 = FSM_dct_8x8_stage_8_0_t81;
    FSM_dct_8x8_stage_8_0_t95[FSM_dct_8x8_stage_8_0_t84 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t94;
    FSM_dct_8x8_stage_8_0_t96 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_8_0_t97 = FSM_dct_8x8_stage_8_0_t96[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t98 = FSM_dct_8x8_stage_8_0_t97[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t99 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_8_0_t100 = FSM_dct_8x8_stage_8_0_t99[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t101 = FSM_dct_8x8_stage_8_0_t100[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t102 = i_data_in[FSM_dct_8x8_stage_8_0_t101 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t103 = FSM_dct_8x8_stage_8_0_t95;
    FSM_dct_8x8_stage_8_0_t103[FSM_dct_8x8_stage_8_0_t98 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t102;
    FSM_dct_8x8_stage_8_0_t104 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_8_0_t105 = FSM_dct_8x8_stage_8_0_t104[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t106 = FSM_dct_8x8_stage_8_0_t105[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t107 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_8_0_t108 = FSM_dct_8x8_stage_8_0_t107[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t109 = FSM_dct_8x8_stage_8_0_t108[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t110 = i_data_in[FSM_dct_8x8_stage_8_0_t109 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t111 = FSM_dct_8x8_stage_8_0_t103;
    FSM_dct_8x8_stage_8_0_t111[FSM_dct_8x8_stage_8_0_t106 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t110;
    FSM_dct_8x8_stage_8_0_t112 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_8_0_t113 = FSM_dct_8x8_stage_8_0_t112[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t114 = FSM_dct_8x8_stage_8_0_t113[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t115 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_8_0_t116 = FSM_dct_8x8_stage_8_0_t115[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t117 = FSM_dct_8x8_stage_8_0_t116[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t118 = i_data_in[FSM_dct_8x8_stage_8_0_t117 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t119 = FSM_dct_8x8_stage_8_0_t111;
    FSM_dct_8x8_stage_8_0_t119[FSM_dct_8x8_stage_8_0_t114 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t118;
    FSM_dct_8x8_stage_8_0_t120 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_8_0_t121 = FSM_dct_8x8_stage_8_0_t120[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t122 = FSM_dct_8x8_stage_8_0_t121[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t123 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_8_0_t124 = FSM_dct_8x8_stage_8_0_t123[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t125 = FSM_dct_8x8_stage_8_0_t124[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t126 = i_data_in[FSM_dct_8x8_stage_8_0_t125 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t127 = FSM_dct_8x8_stage_8_0_t119;
    FSM_dct_8x8_stage_8_0_t127[FSM_dct_8x8_stage_8_0_t122 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t126;
    FSM_dct_8x8_stage_8_0_t128 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_8_0_t129 = FSM_dct_8x8_stage_8_0_t128[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t130 = FSM_dct_8x8_stage_8_0_t129[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t131 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_8_0_t132 = FSM_dct_8x8_stage_8_0_t131[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t133 = FSM_dct_8x8_stage_8_0_t132[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t134 = i_data_in[FSM_dct_8x8_stage_8_0_t133 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t135 = FSM_dct_8x8_stage_8_0_t127;
    FSM_dct_8x8_stage_8_0_t135[FSM_dct_8x8_stage_8_0_t130 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t134;
    FSM_dct_8x8_stage_8_0_t136 = 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_8_0_t137 = FSM_dct_8x8_stage_8_0_t136[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t138 = 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_8_0_t139 = FSM_dct_8x8_stage_8_0_t138[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t140 = i_data_in[FSM_dct_8x8_stage_8_0_t139 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t141 = FSM_dct_8x8_stage_8_0_t135;
    FSM_dct_8x8_stage_8_0_t141[FSM_dct_8x8_stage_8_0_t137 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t140;
    FSM_dct_8x8_stage_8_0_t142 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_8_0_t143 = FSM_dct_8x8_stage_8_0_t142[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t144 = FSM_dct_8x8_stage_8_0_t143[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t145 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_8_0_t146 = FSM_dct_8x8_stage_8_0_t145[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t147 = FSM_dct_8x8_stage_8_0_t146[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t148 = i_data_in[FSM_dct_8x8_stage_8_0_t147 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t149 = FSM_dct_8x8_stage_8_0_t141;
    FSM_dct_8x8_stage_8_0_t149[FSM_dct_8x8_stage_8_0_t144 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t148;
    FSM_dct_8x8_stage_8_0_t150 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_8_0_t151 = FSM_dct_8x8_stage_8_0_t150[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t152 = FSM_dct_8x8_stage_8_0_t151[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t153 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_8_0_t154 = FSM_dct_8x8_stage_8_0_t153[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t155 = FSM_dct_8x8_stage_8_0_t154[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t156 = i_data_in[FSM_dct_8x8_stage_8_0_t155 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t157 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_8_0_t158 = FSM_dct_8x8_stage_8_0_t157[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t159 = FSM_dct_8x8_stage_8_0_t158[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t160 = i_data_in[FSM_dct_8x8_stage_8_0_t159 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t161 = FSM_dct_8x8_stage_8_0_t156 + FSM_dct_8x8_stage_8_0_t160;
    FSM_dct_8x8_stage_8_0_t162 = FSM_dct_8x8_stage_8_0_t161[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t163 = FSM_dct_8x8_stage_8_0_t149;
    FSM_dct_8x8_stage_8_0_t163[FSM_dct_8x8_stage_8_0_t152 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t162;
    FSM_dct_8x8_stage_8_0_t164 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_8_0_t165 = FSM_dct_8x8_stage_8_0_t164[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t166 = FSM_dct_8x8_stage_8_0_t165[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t167 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_8_0_t168 = FSM_dct_8x8_stage_8_0_t167[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t169 = FSM_dct_8x8_stage_8_0_t168[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t170 = i_data_in[FSM_dct_8x8_stage_8_0_t169 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t171 = FSM_dct_8x8_stage_8_0_t163;
    FSM_dct_8x8_stage_8_0_t171[FSM_dct_8x8_stage_8_0_t166 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t170;
    FSM_dct_8x8_stage_8_0_t172 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_8_0_t173 = FSM_dct_8x8_stage_8_0_t172[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t174 = FSM_dct_8x8_stage_8_0_t173[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t175 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_8_0_t176 = FSM_dct_8x8_stage_8_0_t175[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t177 = FSM_dct_8x8_stage_8_0_t176[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t178 = i_data_in[FSM_dct_8x8_stage_8_0_t177 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t179 = FSM_dct_8x8_stage_8_0_t171;
    FSM_dct_8x8_stage_8_0_t179[FSM_dct_8x8_stage_8_0_t174 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t178;
    FSM_dct_8x8_stage_8_0_t180 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_8_0_t181 = FSM_dct_8x8_stage_8_0_t180[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t182 = FSM_dct_8x8_stage_8_0_t181[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t183 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_8_0_t184 = FSM_dct_8x8_stage_8_0_t183[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t185 = FSM_dct_8x8_stage_8_0_t184[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t186 = i_data_in[FSM_dct_8x8_stage_8_0_t185 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t187 = FSM_dct_8x8_stage_8_0_t179;
    FSM_dct_8x8_stage_8_0_t187[FSM_dct_8x8_stage_8_0_t182 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t186;
    FSM_dct_8x8_stage_8_0_t188 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_8_0_t189 = FSM_dct_8x8_stage_8_0_t188[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t190 = FSM_dct_8x8_stage_8_0_t189[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t191 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_8_0_t192 = FSM_dct_8x8_stage_8_0_t191[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t193 = FSM_dct_8x8_stage_8_0_t192[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t194 = i_data_in[FSM_dct_8x8_stage_8_0_t193 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t195 = FSM_dct_8x8_stage_8_0_t187;
    FSM_dct_8x8_stage_8_0_t195[FSM_dct_8x8_stage_8_0_t190 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t194;
    FSM_dct_8x8_stage_8_0_t196 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_8_0_t197 = FSM_dct_8x8_stage_8_0_t196[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t198 = FSM_dct_8x8_stage_8_0_t197[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t199 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_8_0_t200 = FSM_dct_8x8_stage_8_0_t199[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t201 = FSM_dct_8x8_stage_8_0_t200[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t202 = i_data_in[FSM_dct_8x8_stage_8_0_t201 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t203 = FSM_dct_8x8_stage_8_0_t195;
    FSM_dct_8x8_stage_8_0_t203[FSM_dct_8x8_stage_8_0_t198 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t202;
    FSM_dct_8x8_stage_8_0_t204 = 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_8_0_t205 = FSM_dct_8x8_stage_8_0_t204[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t206 = 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_8_0_t207 = FSM_dct_8x8_stage_8_0_t206[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t208 = i_data_in[FSM_dct_8x8_stage_8_0_t207 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t209 = FSM_dct_8x8_stage_8_0_t203;
    FSM_dct_8x8_stage_8_0_t209[FSM_dct_8x8_stage_8_0_t205 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t208;
    FSM_dct_8x8_stage_8_0_t210 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_8_0_t211 = FSM_dct_8x8_stage_8_0_t210[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t212 = FSM_dct_8x8_stage_8_0_t211[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t213 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_8_0_t214 = FSM_dct_8x8_stage_8_0_t213[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t215 = FSM_dct_8x8_stage_8_0_t214[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t216 = i_data_in[FSM_dct_8x8_stage_8_0_t215 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t217 = FSM_dct_8x8_stage_8_0_t209;
    FSM_dct_8x8_stage_8_0_t217[FSM_dct_8x8_stage_8_0_t212 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t216;
    FSM_dct_8x8_stage_8_0_t218 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_8_0_t219 = FSM_dct_8x8_stage_8_0_t218[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t220 = FSM_dct_8x8_stage_8_0_t219[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t221 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_8_0_t222 = FSM_dct_8x8_stage_8_0_t221[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t223 = FSM_dct_8x8_stage_8_0_t222[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t224 = i_data_in[FSM_dct_8x8_stage_8_0_t223 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t225 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_8_0_t226 = FSM_dct_8x8_stage_8_0_t225[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t227 = FSM_dct_8x8_stage_8_0_t226[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t228 = i_data_in[FSM_dct_8x8_stage_8_0_t227 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t229 = FSM_dct_8x8_stage_8_0_t224 + FSM_dct_8x8_stage_8_0_t228;
    FSM_dct_8x8_stage_8_0_t230 = FSM_dct_8x8_stage_8_0_t229[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t231 = FSM_dct_8x8_stage_8_0_t217;
    FSM_dct_8x8_stage_8_0_t231[FSM_dct_8x8_stage_8_0_t220 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t230;
    FSM_dct_8x8_stage_8_0_t232 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_8_0_t233 = FSM_dct_8x8_stage_8_0_t232[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t234 = FSM_dct_8x8_stage_8_0_t233[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t235 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_8_0_t236 = FSM_dct_8x8_stage_8_0_t235[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t237 = FSM_dct_8x8_stage_8_0_t236[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t238 = i_data_in[FSM_dct_8x8_stage_8_0_t237 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t239 = FSM_dct_8x8_stage_8_0_t231;
    FSM_dct_8x8_stage_8_0_t239[FSM_dct_8x8_stage_8_0_t234 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t238;
    FSM_dct_8x8_stage_8_0_t240 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_8_0_t241 = FSM_dct_8x8_stage_8_0_t240[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t242 = FSM_dct_8x8_stage_8_0_t241[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t243 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_8_0_t244 = FSM_dct_8x8_stage_8_0_t243[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t245 = FSM_dct_8x8_stage_8_0_t244[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t246 = i_data_in[FSM_dct_8x8_stage_8_0_t245 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t247 = FSM_dct_8x8_stage_8_0_t239;
    FSM_dct_8x8_stage_8_0_t247[FSM_dct_8x8_stage_8_0_t242 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t246;
    FSM_dct_8x8_stage_8_0_t248 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_8_0_t249 = FSM_dct_8x8_stage_8_0_t248[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t250 = FSM_dct_8x8_stage_8_0_t249[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t251 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_8_0_t252 = FSM_dct_8x8_stage_8_0_t251[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t253 = FSM_dct_8x8_stage_8_0_t252[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t254 = i_data_in[FSM_dct_8x8_stage_8_0_t253 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t255 = FSM_dct_8x8_stage_8_0_t247;
    FSM_dct_8x8_stage_8_0_t255[FSM_dct_8x8_stage_8_0_t250 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t254;
    FSM_dct_8x8_stage_8_0_t256 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_8_0_t257 = FSM_dct_8x8_stage_8_0_t256[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t258 = FSM_dct_8x8_stage_8_0_t257[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t259 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_8_0_t260 = FSM_dct_8x8_stage_8_0_t259[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t261 = FSM_dct_8x8_stage_8_0_t260[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t262 = i_data_in[FSM_dct_8x8_stage_8_0_t261 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t263 = FSM_dct_8x8_stage_8_0_t255;
    FSM_dct_8x8_stage_8_0_t263[FSM_dct_8x8_stage_8_0_t258 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t262;
    FSM_dct_8x8_stage_8_0_t264 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_8_0_t265 = FSM_dct_8x8_stage_8_0_t264[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t266 = FSM_dct_8x8_stage_8_0_t265[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t267 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_8_0_t268 = FSM_dct_8x8_stage_8_0_t267[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t269 = FSM_dct_8x8_stage_8_0_t268[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t270 = i_data_in[FSM_dct_8x8_stage_8_0_t269 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t271 = FSM_dct_8x8_stage_8_0_t263;
    FSM_dct_8x8_stage_8_0_t271[FSM_dct_8x8_stage_8_0_t266 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t270;
    FSM_dct_8x8_stage_8_0_t272 = 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_8_0_t273 = FSM_dct_8x8_stage_8_0_t272[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t274 = 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_8_0_t275 = FSM_dct_8x8_stage_8_0_t274[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t276 = i_data_in[FSM_dct_8x8_stage_8_0_t275 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t277 = FSM_dct_8x8_stage_8_0_t271;
    FSM_dct_8x8_stage_8_0_t277[FSM_dct_8x8_stage_8_0_t273 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t276;
    FSM_dct_8x8_stage_8_0_t278 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_8_0_t279 = FSM_dct_8x8_stage_8_0_t278[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t280 = FSM_dct_8x8_stage_8_0_t279[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t281 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_8_0_t282 = FSM_dct_8x8_stage_8_0_t281[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t283 = FSM_dct_8x8_stage_8_0_t282[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t284 = i_data_in[FSM_dct_8x8_stage_8_0_t283 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t285 = FSM_dct_8x8_stage_8_0_t277;
    FSM_dct_8x8_stage_8_0_t285[FSM_dct_8x8_stage_8_0_t280 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t284;
    FSM_dct_8x8_stage_8_0_t286 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_8_0_t287 = FSM_dct_8x8_stage_8_0_t286[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t288 = FSM_dct_8x8_stage_8_0_t287[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t289 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_8_0_t290 = FSM_dct_8x8_stage_8_0_t289[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t291 = FSM_dct_8x8_stage_8_0_t290[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t292 = i_data_in[FSM_dct_8x8_stage_8_0_t291 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t293 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_8_0_t294 = FSM_dct_8x8_stage_8_0_t293[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t295 = FSM_dct_8x8_stage_8_0_t294[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t296 = i_data_in[FSM_dct_8x8_stage_8_0_t295 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t297 = FSM_dct_8x8_stage_8_0_t292 + FSM_dct_8x8_stage_8_0_t296;
    FSM_dct_8x8_stage_8_0_t298 = FSM_dct_8x8_stage_8_0_t297[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t299 = FSM_dct_8x8_stage_8_0_t285;
    FSM_dct_8x8_stage_8_0_t299[FSM_dct_8x8_stage_8_0_t288 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t298;
    FSM_dct_8x8_stage_8_0_t300 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_8_0_t301 = FSM_dct_8x8_stage_8_0_t300[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t302 = FSM_dct_8x8_stage_8_0_t301[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t303 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_8_0_t304 = FSM_dct_8x8_stage_8_0_t303[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t305 = FSM_dct_8x8_stage_8_0_t304[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t306 = i_data_in[FSM_dct_8x8_stage_8_0_t305 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t307 = FSM_dct_8x8_stage_8_0_t299;
    FSM_dct_8x8_stage_8_0_t307[FSM_dct_8x8_stage_8_0_t302 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t306;
    FSM_dct_8x8_stage_8_0_t308 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_8_0_t309 = FSM_dct_8x8_stage_8_0_t308[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t310 = FSM_dct_8x8_stage_8_0_t309[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t311 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_8_0_t312 = FSM_dct_8x8_stage_8_0_t311[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t313 = FSM_dct_8x8_stage_8_0_t312[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t314 = i_data_in[FSM_dct_8x8_stage_8_0_t313 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t315 = FSM_dct_8x8_stage_8_0_t307;
    FSM_dct_8x8_stage_8_0_t315[FSM_dct_8x8_stage_8_0_t310 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t314;
    FSM_dct_8x8_stage_8_0_t316 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_8_0_t317 = FSM_dct_8x8_stage_8_0_t316[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t318 = FSM_dct_8x8_stage_8_0_t317[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t319 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_8_0_t320 = FSM_dct_8x8_stage_8_0_t319[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t321 = FSM_dct_8x8_stage_8_0_t320[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t322 = i_data_in[FSM_dct_8x8_stage_8_0_t321 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t323 = FSM_dct_8x8_stage_8_0_t315;
    FSM_dct_8x8_stage_8_0_t323[FSM_dct_8x8_stage_8_0_t318 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t322;
    FSM_dct_8x8_stage_8_0_t324 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_8_0_t325 = FSM_dct_8x8_stage_8_0_t324[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t326 = FSM_dct_8x8_stage_8_0_t325[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t327 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_8_0_t328 = FSM_dct_8x8_stage_8_0_t327[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t329 = FSM_dct_8x8_stage_8_0_t328[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t330 = i_data_in[FSM_dct_8x8_stage_8_0_t329 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t331 = FSM_dct_8x8_stage_8_0_t323;
    FSM_dct_8x8_stage_8_0_t331[FSM_dct_8x8_stage_8_0_t326 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t330;
    FSM_dct_8x8_stage_8_0_t332 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_8_0_t333 = FSM_dct_8x8_stage_8_0_t332[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t334 = FSM_dct_8x8_stage_8_0_t333[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t335 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_8_0_t336 = FSM_dct_8x8_stage_8_0_t335[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t337 = FSM_dct_8x8_stage_8_0_t336[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t338 = i_data_in[FSM_dct_8x8_stage_8_0_t337 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t339 = FSM_dct_8x8_stage_8_0_t331;
    FSM_dct_8x8_stage_8_0_t339[FSM_dct_8x8_stage_8_0_t334 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t338;
    FSM_dct_8x8_stage_8_0_t340 = 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_8_0_t341 = FSM_dct_8x8_stage_8_0_t340[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t342 = 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_8_0_t343 = FSM_dct_8x8_stage_8_0_t342[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t344 = i_data_in[FSM_dct_8x8_stage_8_0_t343 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t345 = FSM_dct_8x8_stage_8_0_t339;
    FSM_dct_8x8_stage_8_0_t345[FSM_dct_8x8_stage_8_0_t341 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t344;
    FSM_dct_8x8_stage_8_0_t346 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_8_0_t347 = FSM_dct_8x8_stage_8_0_t346[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t348 = FSM_dct_8x8_stage_8_0_t347[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t349 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_8_0_t350 = FSM_dct_8x8_stage_8_0_t349[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t351 = FSM_dct_8x8_stage_8_0_t350[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t352 = i_data_in[FSM_dct_8x8_stage_8_0_t351 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t353 = FSM_dct_8x8_stage_8_0_t345;
    FSM_dct_8x8_stage_8_0_t353[FSM_dct_8x8_stage_8_0_t348 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t352;
    FSM_dct_8x8_stage_8_0_t354 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_8_0_t355 = FSM_dct_8x8_stage_8_0_t354[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t356 = FSM_dct_8x8_stage_8_0_t355[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t357 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_8_0_t358 = FSM_dct_8x8_stage_8_0_t357[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t359 = FSM_dct_8x8_stage_8_0_t358[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t360 = i_data_in[FSM_dct_8x8_stage_8_0_t359 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t361 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_8_0_t362 = FSM_dct_8x8_stage_8_0_t361[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t363 = FSM_dct_8x8_stage_8_0_t362[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t364 = i_data_in[FSM_dct_8x8_stage_8_0_t363 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t365 = FSM_dct_8x8_stage_8_0_t360 + FSM_dct_8x8_stage_8_0_t364;
    FSM_dct_8x8_stage_8_0_t366 = FSM_dct_8x8_stage_8_0_t365[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t367 = FSM_dct_8x8_stage_8_0_t353;
    FSM_dct_8x8_stage_8_0_t367[FSM_dct_8x8_stage_8_0_t356 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t366;
    FSM_dct_8x8_stage_8_0_t368 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_8_0_t369 = FSM_dct_8x8_stage_8_0_t368[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t370 = FSM_dct_8x8_stage_8_0_t369[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t371 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_8_0_t372 = FSM_dct_8x8_stage_8_0_t371[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t373 = FSM_dct_8x8_stage_8_0_t372[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t374 = i_data_in[FSM_dct_8x8_stage_8_0_t373 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t375 = FSM_dct_8x8_stage_8_0_t367;
    FSM_dct_8x8_stage_8_0_t375[FSM_dct_8x8_stage_8_0_t370 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t374;
    FSM_dct_8x8_stage_8_0_t376 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_8_0_t377 = FSM_dct_8x8_stage_8_0_t376[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t378 = FSM_dct_8x8_stage_8_0_t377[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t379 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_8_0_t380 = FSM_dct_8x8_stage_8_0_t379[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t381 = FSM_dct_8x8_stage_8_0_t380[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t382 = i_data_in[FSM_dct_8x8_stage_8_0_t381 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t383 = FSM_dct_8x8_stage_8_0_t375;
    FSM_dct_8x8_stage_8_0_t383[FSM_dct_8x8_stage_8_0_t378 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t382;
    FSM_dct_8x8_stage_8_0_t384 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_8_0_t385 = FSM_dct_8x8_stage_8_0_t384[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t386 = FSM_dct_8x8_stage_8_0_t385[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t387 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_8_0_t388 = FSM_dct_8x8_stage_8_0_t387[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t389 = FSM_dct_8x8_stage_8_0_t388[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t390 = i_data_in[FSM_dct_8x8_stage_8_0_t389 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t391 = FSM_dct_8x8_stage_8_0_t383;
    FSM_dct_8x8_stage_8_0_t391[FSM_dct_8x8_stage_8_0_t386 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t390;
    FSM_dct_8x8_stage_8_0_t392 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_8_0_t393 = FSM_dct_8x8_stage_8_0_t392[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t394 = FSM_dct_8x8_stage_8_0_t393[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t395 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_8_0_t396 = FSM_dct_8x8_stage_8_0_t395[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t397 = FSM_dct_8x8_stage_8_0_t396[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t398 = i_data_in[FSM_dct_8x8_stage_8_0_t397 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t399 = FSM_dct_8x8_stage_8_0_t391;
    FSM_dct_8x8_stage_8_0_t399[FSM_dct_8x8_stage_8_0_t394 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t398;
    FSM_dct_8x8_stage_8_0_t400 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_8_0_t401 = FSM_dct_8x8_stage_8_0_t400[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t402 = FSM_dct_8x8_stage_8_0_t401[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t403 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_8_0_t404 = FSM_dct_8x8_stage_8_0_t403[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t405 = FSM_dct_8x8_stage_8_0_t404[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t406 = i_data_in[FSM_dct_8x8_stage_8_0_t405 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t407 = FSM_dct_8x8_stage_8_0_t399;
    FSM_dct_8x8_stage_8_0_t407[FSM_dct_8x8_stage_8_0_t402 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t406;
    FSM_dct_8x8_stage_8_0_t408 = 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_8_0_t409 = FSM_dct_8x8_stage_8_0_t408[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t410 = 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_8_0_t411 = FSM_dct_8x8_stage_8_0_t410[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t412 = i_data_in[FSM_dct_8x8_stage_8_0_t411 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t413 = FSM_dct_8x8_stage_8_0_t407;
    FSM_dct_8x8_stage_8_0_t413[FSM_dct_8x8_stage_8_0_t409 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t412;
    FSM_dct_8x8_stage_8_0_t414 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_8_0_t415 = FSM_dct_8x8_stage_8_0_t414[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t416 = FSM_dct_8x8_stage_8_0_t415[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t417 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_8_0_t418 = FSM_dct_8x8_stage_8_0_t417[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t419 = FSM_dct_8x8_stage_8_0_t418[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t420 = i_data_in[FSM_dct_8x8_stage_8_0_t419 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t421 = FSM_dct_8x8_stage_8_0_t413;
    FSM_dct_8x8_stage_8_0_t421[FSM_dct_8x8_stage_8_0_t416 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t420;
    FSM_dct_8x8_stage_8_0_t422 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_8_0_t423 = FSM_dct_8x8_stage_8_0_t422[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t424 = FSM_dct_8x8_stage_8_0_t423[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t425 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_8_0_t426 = FSM_dct_8x8_stage_8_0_t425[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t427 = FSM_dct_8x8_stage_8_0_t426[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t428 = i_data_in[FSM_dct_8x8_stage_8_0_t427 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t429 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_8_0_t430 = FSM_dct_8x8_stage_8_0_t429[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t431 = FSM_dct_8x8_stage_8_0_t430[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t432 = i_data_in[FSM_dct_8x8_stage_8_0_t431 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t433 = FSM_dct_8x8_stage_8_0_t428 + FSM_dct_8x8_stage_8_0_t432;
    FSM_dct_8x8_stage_8_0_t434 = FSM_dct_8x8_stage_8_0_t433[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t435 = FSM_dct_8x8_stage_8_0_t421;
    FSM_dct_8x8_stage_8_0_t435[FSM_dct_8x8_stage_8_0_t424 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t434;
    FSM_dct_8x8_stage_8_0_t436 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_8_0_t437 = FSM_dct_8x8_stage_8_0_t436[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t438 = FSM_dct_8x8_stage_8_0_t437[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t439 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_8_0_t440 = FSM_dct_8x8_stage_8_0_t439[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t441 = FSM_dct_8x8_stage_8_0_t440[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t442 = i_data_in[FSM_dct_8x8_stage_8_0_t441 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t443 = FSM_dct_8x8_stage_8_0_t435;
    FSM_dct_8x8_stage_8_0_t443[FSM_dct_8x8_stage_8_0_t438 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t442;
    FSM_dct_8x8_stage_8_0_t444 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_8_0_t445 = FSM_dct_8x8_stage_8_0_t444[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t446 = FSM_dct_8x8_stage_8_0_t445[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t447 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_8_0_t448 = FSM_dct_8x8_stage_8_0_t447[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t449 = FSM_dct_8x8_stage_8_0_t448[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t450 = i_data_in[FSM_dct_8x8_stage_8_0_t449 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t451 = FSM_dct_8x8_stage_8_0_t443;
    FSM_dct_8x8_stage_8_0_t451[FSM_dct_8x8_stage_8_0_t446 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t450;
    FSM_dct_8x8_stage_8_0_t452 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_8_0_t453 = FSM_dct_8x8_stage_8_0_t452[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t454 = FSM_dct_8x8_stage_8_0_t453[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t455 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_8_0_t456 = FSM_dct_8x8_stage_8_0_t455[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t457 = FSM_dct_8x8_stage_8_0_t456[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t458 = i_data_in[FSM_dct_8x8_stage_8_0_t457 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t459 = FSM_dct_8x8_stage_8_0_t451;
    FSM_dct_8x8_stage_8_0_t459[FSM_dct_8x8_stage_8_0_t454 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t458;
    FSM_dct_8x8_stage_8_0_t460 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_8_0_t461 = FSM_dct_8x8_stage_8_0_t460[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t462 = FSM_dct_8x8_stage_8_0_t461[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t463 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_8_0_t464 = FSM_dct_8x8_stage_8_0_t463[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t465 = FSM_dct_8x8_stage_8_0_t464[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t466 = i_data_in[FSM_dct_8x8_stage_8_0_t465 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t467 = FSM_dct_8x8_stage_8_0_t459;
    FSM_dct_8x8_stage_8_0_t467[FSM_dct_8x8_stage_8_0_t462 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t466;
    FSM_dct_8x8_stage_8_0_t468 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_8_0_t469 = FSM_dct_8x8_stage_8_0_t468[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t470 = FSM_dct_8x8_stage_8_0_t469[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t471 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_8_0_t472 = FSM_dct_8x8_stage_8_0_t471[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t473 = FSM_dct_8x8_stage_8_0_t472[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t474 = i_data_in[FSM_dct_8x8_stage_8_0_t473 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t475 = FSM_dct_8x8_stage_8_0_t467;
    FSM_dct_8x8_stage_8_0_t475[FSM_dct_8x8_stage_8_0_t470 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t474;
    FSM_dct_8x8_stage_8_0_t476 = 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_8_0_t477 = FSM_dct_8x8_stage_8_0_t476[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t478 = 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_8_0_t479 = FSM_dct_8x8_stage_8_0_t478[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t480 = i_data_in[FSM_dct_8x8_stage_8_0_t479 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t481 = FSM_dct_8x8_stage_8_0_t475;
    FSM_dct_8x8_stage_8_0_t481[FSM_dct_8x8_stage_8_0_t477 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t480;
    FSM_dct_8x8_stage_8_0_t482 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_8_0_t483 = FSM_dct_8x8_stage_8_0_t482[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t484 = FSM_dct_8x8_stage_8_0_t483[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t485 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_8_0_t486 = FSM_dct_8x8_stage_8_0_t485[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t487 = FSM_dct_8x8_stage_8_0_t486[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t488 = i_data_in[FSM_dct_8x8_stage_8_0_t487 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t489 = FSM_dct_8x8_stage_8_0_t481;
    FSM_dct_8x8_stage_8_0_t489[FSM_dct_8x8_stage_8_0_t484 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t488;
    FSM_dct_8x8_stage_8_0_t490 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_8_0_t491 = FSM_dct_8x8_stage_8_0_t490[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t492 = FSM_dct_8x8_stage_8_0_t491[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t493 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_8_0_t494 = FSM_dct_8x8_stage_8_0_t493[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t495 = FSM_dct_8x8_stage_8_0_t494[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t496 = i_data_in[FSM_dct_8x8_stage_8_0_t495 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t497 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_8_0_t498 = FSM_dct_8x8_stage_8_0_t497[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t499 = FSM_dct_8x8_stage_8_0_t498[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t500 = i_data_in[FSM_dct_8x8_stage_8_0_t499 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t501 = FSM_dct_8x8_stage_8_0_t496 + FSM_dct_8x8_stage_8_0_t500;
    FSM_dct_8x8_stage_8_0_t502 = FSM_dct_8x8_stage_8_0_t501[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t503 = FSM_dct_8x8_stage_8_0_t489;
    FSM_dct_8x8_stage_8_0_t503[FSM_dct_8x8_stage_8_0_t492 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t502;
    FSM_dct_8x8_stage_8_0_t504 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_8_0_t505 = FSM_dct_8x8_stage_8_0_t504[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t506 = FSM_dct_8x8_stage_8_0_t505[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t507 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_8_0_t508 = FSM_dct_8x8_stage_8_0_t507[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t509 = FSM_dct_8x8_stage_8_0_t508[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t510 = i_data_in[FSM_dct_8x8_stage_8_0_t509 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t511 = FSM_dct_8x8_stage_8_0_t503;
    FSM_dct_8x8_stage_8_0_t511[FSM_dct_8x8_stage_8_0_t506 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t510;
    FSM_dct_8x8_stage_8_0_t512 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_8_0_t513 = FSM_dct_8x8_stage_8_0_t512[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t514 = FSM_dct_8x8_stage_8_0_t513[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t515 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_8_0_t516 = FSM_dct_8x8_stage_8_0_t515[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t517 = FSM_dct_8x8_stage_8_0_t516[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t518 = i_data_in[FSM_dct_8x8_stage_8_0_t517 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t519 = FSM_dct_8x8_stage_8_0_t511;
    FSM_dct_8x8_stage_8_0_t519[FSM_dct_8x8_stage_8_0_t514 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t518;
    FSM_dct_8x8_stage_8_0_t520 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_8_0_t521 = FSM_dct_8x8_stage_8_0_t520[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t522 = FSM_dct_8x8_stage_8_0_t521[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t523 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_8_0_t524 = FSM_dct_8x8_stage_8_0_t523[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t525 = FSM_dct_8x8_stage_8_0_t524[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t526 = i_data_in[FSM_dct_8x8_stage_8_0_t525 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t527 = FSM_dct_8x8_stage_8_0_t519;
    FSM_dct_8x8_stage_8_0_t527[FSM_dct_8x8_stage_8_0_t522 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t526;
    FSM_dct_8x8_stage_8_0_t528 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_8_0_t529 = FSM_dct_8x8_stage_8_0_t528[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t530 = FSM_dct_8x8_stage_8_0_t529[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t531 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_8_0_t532 = FSM_dct_8x8_stage_8_0_t531[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t533 = FSM_dct_8x8_stage_8_0_t532[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t534 = i_data_in[FSM_dct_8x8_stage_8_0_t533 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t535 = FSM_dct_8x8_stage_8_0_t527;
    FSM_dct_8x8_stage_8_0_t535[FSM_dct_8x8_stage_8_0_t530 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t534;
    FSM_dct_8x8_stage_8_0_t536 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_8_0_t537 = FSM_dct_8x8_stage_8_0_t536[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t538 = FSM_dct_8x8_stage_8_0_t537[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t539 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_8_0_t540 = FSM_dct_8x8_stage_8_0_t539[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_8_0_t541 = FSM_dct_8x8_stage_8_0_t540[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_8_0_t542 = i_data_in[FSM_dct_8x8_stage_8_0_t541 * 32 +: 32];
    FSM_dct_8x8_stage_8_0_t543 = FSM_dct_8x8_stage_8_0_t535;
    FSM_dct_8x8_stage_8_0_t543[FSM_dct_8x8_stage_8_0_t538 * 32 +: 32] = FSM_dct_8x8_stage_8_0_t542;
end

assign FSM_dct_8x8_stage_8_0_in_ready = 1'b1;

always @(posedge clk) begin
    FSM_dct_8x8_stage_8_0_st_dummy_reg <= FSM_dct_8x8_stage_8_0_st_dummy_reg;
    if (rst) begin
        FSM_dct_8x8_stage_8_0_st_dummy_reg <= 32'b0;
    end
end
/* End submodules of dct_8x8_stage_8 */
/* End module dct_8x8_stage_8 */
endgenerate
endmodule
