`timescale 1ns / 1ps

module shift_rows_inner
(
    input wire clk,
    input wire rst,
    input wire [64-1:0] i_higher_bits,
    input wire [64-1:0] i_lower_bits,
    input wire i_valid,
    output wire i_ready,
    output wire [64-1:0] o_data_out_higher,
    output wire [64-1:0] o_data_out_lower,
    output wire o_valid,
    input wire o_ready
);

generate
/*
    Begin module shift_rows
*/
/*
    Wires declared by shift_rows
*/
wire FSM_shift_rows_0_in_ready;
wire [64-1:0] FSM_shift_rows_0_out_data_out_higher;
wire [64-1:0] FSM_shift_rows_0_out_data_out_lower;
wire FSM_shift_rows_0_out_valid;
/* End wires declared by shift_rows */

/*
    Wiring by shift_rows
*/
assign i_ready = FSM_shift_rows_0_in_ready;
assign o_data_out_higher = FSM_shift_rows_0_out_data_out_higher;
assign o_data_out_lower = FSM_shift_rows_0_out_data_out_lower;
assign o_valid = FSM_shift_rows_0_out_valid;
/* End wiring by shift_rows */

/*
    Submodules of shift_rows
*/
reg [64-1:0] FSM_shift_rows_0_st_dummy_reg = 64'b0;

reg [1024-1:0] FSM_shift_rows_0_t0;
reg [64-1:0] FSM_shift_rows_0_t1;
reg [6-1:0] FSM_shift_rows_0_t2;
reg [64-1:0] FSM_shift_rows_0_t3;
reg [6-1:0] FSM_shift_rows_0_t4;
reg [64-1:0] FSM_shift_rows_0_t5;
reg [6-1:0] FSM_shift_rows_0_t6;
reg [64-1:0] FSM_shift_rows_0_t7;
reg [6-1:0] FSM_shift_rows_0_t8;
reg [64-1:0] FSM_shift_rows_0_t9;
reg [6-1:0] FSM_shift_rows_0_t10;
reg [64-1:0] FSM_shift_rows_0_t11;
reg [6-1:0] FSM_shift_rows_0_t12;
reg [64-1:0] FSM_shift_rows_0_t13;
reg [6-1:0] FSM_shift_rows_0_t14;
reg [64-1:0] FSM_shift_rows_0_t15;
reg [6-1:0] FSM_shift_rows_0_t16;
reg [64-1:0] FSM_shift_rows_0_t17;
reg [6-1:0] FSM_shift_rows_0_t18;
reg [64-1:0] FSM_shift_rows_0_t19;
reg [6-1:0] FSM_shift_rows_0_t20;
reg [64-1:0] FSM_shift_rows_0_t21;
reg [6-1:0] FSM_shift_rows_0_t22;
reg [64-1:0] FSM_shift_rows_0_t23;
reg [6-1:0] FSM_shift_rows_0_t24;
reg [64-1:0] FSM_shift_rows_0_t25;
reg [6-1:0] FSM_shift_rows_0_t26;
reg [64-1:0] FSM_shift_rows_0_t27;
reg [6-1:0] FSM_shift_rows_0_t28;
reg [64-1:0] FSM_shift_rows_0_t29;
reg [4-1:0] FSM_shift_rows_0_t30;
reg [64-1:0] FSM_shift_rows_0_t31;
reg [64-1:0] FSM_shift_rows_0_t32;
reg [6-1:0] FSM_shift_rows_0_t33;
reg [64-1:0] FSM_shift_rows_0_t34;
reg [4-1:0] FSM_shift_rows_0_t35;
reg [64-1:0] FSM_shift_rows_0_t36;
reg [64-1:0] FSM_shift_rows_0_t37;
reg [6-1:0] FSM_shift_rows_0_t38;
reg [64-1:0] FSM_shift_rows_0_t39;
reg [4-1:0] FSM_shift_rows_0_t40;
reg [64-1:0] FSM_shift_rows_0_t41;
reg [64-1:0] FSM_shift_rows_0_t42;
reg [6-1:0] FSM_shift_rows_0_t43;
reg [64-1:0] FSM_shift_rows_0_t44;
reg [4-1:0] FSM_shift_rows_0_t45;
reg [64-1:0] FSM_shift_rows_0_t46;
reg [64-1:0] FSM_shift_rows_0_t47;
reg [6-1:0] FSM_shift_rows_0_t48;
reg [64-1:0] FSM_shift_rows_0_t49;
reg [4-1:0] FSM_shift_rows_0_t50;
reg [64-1:0] FSM_shift_rows_0_t51;
reg [64-1:0] FSM_shift_rows_0_t52;
reg [6-1:0] FSM_shift_rows_0_t53;
reg [64-1:0] FSM_shift_rows_0_t54;
reg [4-1:0] FSM_shift_rows_0_t55;
reg [64-1:0] FSM_shift_rows_0_t56;
reg [64-1:0] FSM_shift_rows_0_t57;
reg [6-1:0] FSM_shift_rows_0_t58;
reg [64-1:0] FSM_shift_rows_0_t59;
reg [4-1:0] FSM_shift_rows_0_t60;
reg [64-1:0] FSM_shift_rows_0_t61;
reg [64-1:0] FSM_shift_rows_0_t62;
reg [6-1:0] FSM_shift_rows_0_t63;
reg [64-1:0] FSM_shift_rows_0_t64;
reg [4-1:0] FSM_shift_rows_0_t65;
reg [64-1:0] FSM_shift_rows_0_t66;
reg [64-1:0] FSM_shift_rows_0_t67;
reg [4-1:0] FSM_shift_rows_0_t68;
reg [64-1:0] FSM_shift_rows_0_t69;
reg [64-1:0] FSM_shift_rows_0_t70;
reg [6-1:0] FSM_shift_rows_0_t71;
reg [64-1:0] FSM_shift_rows_0_t72;
reg [4-1:0] FSM_shift_rows_0_t73;
reg [64-1:0] FSM_shift_rows_0_t74;
reg [64-1:0] FSM_shift_rows_0_t75;
reg [6-1:0] FSM_shift_rows_0_t76;
reg [64-1:0] FSM_shift_rows_0_t77;
reg [4-1:0] FSM_shift_rows_0_t78;
reg [64-1:0] FSM_shift_rows_0_t79;
reg [64-1:0] FSM_shift_rows_0_t80;
reg [6-1:0] FSM_shift_rows_0_t81;
reg [64-1:0] FSM_shift_rows_0_t82;
reg [4-1:0] FSM_shift_rows_0_t83;
reg [64-1:0] FSM_shift_rows_0_t84;
reg [64-1:0] FSM_shift_rows_0_t85;
reg [6-1:0] FSM_shift_rows_0_t86;
reg [64-1:0] FSM_shift_rows_0_t87;
reg [4-1:0] FSM_shift_rows_0_t88;
reg [64-1:0] FSM_shift_rows_0_t89;
reg [64-1:0] FSM_shift_rows_0_t90;
reg [6-1:0] FSM_shift_rows_0_t91;
reg [64-1:0] FSM_shift_rows_0_t92;
reg [4-1:0] FSM_shift_rows_0_t93;
reg [64-1:0] FSM_shift_rows_0_t94;
reg [64-1:0] FSM_shift_rows_0_t95;
reg [6-1:0] FSM_shift_rows_0_t96;
reg [64-1:0] FSM_shift_rows_0_t97;
reg [4-1:0] FSM_shift_rows_0_t98;
reg [64-1:0] FSM_shift_rows_0_t99;
reg [64-1:0] FSM_shift_rows_0_t100;
reg [6-1:0] FSM_shift_rows_0_t101;
reg [64-1:0] FSM_shift_rows_0_t102;
reg [4-1:0] FSM_shift_rows_0_t103;
reg [64-1:0] FSM_shift_rows_0_t104;

assign FSM_shift_rows_0_out_data_out_higher = (FSM_shift_rows_0_t31 << FSM_shift_rows_0_t33) | ((FSM_shift_rows_0_t36 << FSM_shift_rows_0_t38) | ((FSM_shift_rows_0_t41 << FSM_shift_rows_0_t43) | ((FSM_shift_rows_0_t46 << FSM_shift_rows_0_t48) | ((FSM_shift_rows_0_t51 << FSM_shift_rows_0_t53) | ((FSM_shift_rows_0_t56 << FSM_shift_rows_0_t58) | ((FSM_shift_rows_0_t61 << FSM_shift_rows_0_t63) | FSM_shift_rows_0_t66))))));
assign FSM_shift_rows_0_out_data_out_lower = (FSM_shift_rows_0_t69 << FSM_shift_rows_0_t71) | ((FSM_shift_rows_0_t74 << FSM_shift_rows_0_t76) | ((FSM_shift_rows_0_t79 << FSM_shift_rows_0_t81) | ((FSM_shift_rows_0_t84 << FSM_shift_rows_0_t86) | ((FSM_shift_rows_0_t89 << FSM_shift_rows_0_t91) | ((FSM_shift_rows_0_t94 << FSM_shift_rows_0_t96) | ((FSM_shift_rows_0_t99 << FSM_shift_rows_0_t101) | FSM_shift_rows_0_t104))))));
assign FSM_shift_rows_0_out_valid = 1'b1;

initial begin
    FSM_shift_rows_0_t0[0 * 64 +: 64] = i_lower_bits & 64'b0000000000000000000000000000000000000000000000000000000011111111;
    FSM_shift_rows_0_t1 = 64'b0000000000000000000000000000000000000000000000000000000000001000;
    FSM_shift_rows_0_t2 = FSM_shift_rows_0_t1[6'b0 * 1 +: 6 * 1];
    FSM_shift_rows_0_t0[1 * 64 +: 64] = (i_lower_bits >> FSM_shift_rows_0_t2) & 64'b0000000000000000000000000000000000000000000000000000000011111111;
    FSM_shift_rows_0_t3 = 64'b0000000000000000000000000000000000000000000000000000000000010000;
    FSM_shift_rows_0_t4 = FSM_shift_rows_0_t3[6'b0 * 1 +: 6 * 1];
    FSM_shift_rows_0_t0[2 * 64 +: 64] = (i_lower_bits >> FSM_shift_rows_0_t4) & 64'b0000000000000000000000000000000000000000000000000000000011111111;
    FSM_shift_rows_0_t5 = 64'b0000000000000000000000000000000000000000000000000000000000011000;
    FSM_shift_rows_0_t6 = FSM_shift_rows_0_t5[6'b0 * 1 +: 6 * 1];
    FSM_shift_rows_0_t0[3 * 64 +: 64] = (i_lower_bits >> FSM_shift_rows_0_t6) & 64'b0000000000000000000000000000000000000000000000000000000011111111;
    FSM_shift_rows_0_t7 = 64'b0000000000000000000000000000000000000000000000000000000000101000;
    FSM_shift_rows_0_t8 = FSM_shift_rows_0_t7[6'b0 * 1 +: 6 * 1];
    FSM_shift_rows_0_t0[4 * 64 +: 64] = (i_lower_bits >> FSM_shift_rows_0_t8) & 64'b0000000000000000000000000000000000000000000000000000000011111111;
    FSM_shift_rows_0_t9 = 64'b0000000000000000000000000000000000000000000000000000000000110000;
    FSM_shift_rows_0_t10 = FSM_shift_rows_0_t9[6'b0 * 1 +: 6 * 1];
    FSM_shift_rows_0_t0[5 * 64 +: 64] = (i_lower_bits >> FSM_shift_rows_0_t10) & 64'b0000000000000000000000000000000000000000000000000000000011111111;
    FSM_shift_rows_0_t11 = 64'b0000000000000000000000000000000000000000000000000000000000111000;
    FSM_shift_rows_0_t12 = FSM_shift_rows_0_t11[6'b0 * 1 +: 6 * 1];
    FSM_shift_rows_0_t0[6 * 64 +: 64] = (i_lower_bits >> FSM_shift_rows_0_t12) & 64'b0000000000000000000000000000000000000000000000000000000011111111;
    FSM_shift_rows_0_t13 = 64'b0000000000000000000000000000000000000000000000000000000000100000;
    FSM_shift_rows_0_t14 = FSM_shift_rows_0_t13[6'b0 * 1 +: 6 * 1];
    FSM_shift_rows_0_t0[7 * 64 +: 64] = (i_lower_bits >> FSM_shift_rows_0_t14) & 64'b0000000000000000000000000000000000000000000000000000000011111111;
    FSM_shift_rows_0_t15 = 64'b0000000000000000000000000000000000000000000000000000000000010000;
    FSM_shift_rows_0_t16 = FSM_shift_rows_0_t15[6'b0 * 1 +: 6 * 1];
    FSM_shift_rows_0_t0[8 * 64 +: 64] = (i_higher_bits >> FSM_shift_rows_0_t16) & 64'b0000000000000000000000000000000000000000000000000000000011111111;
    FSM_shift_rows_0_t17 = 64'b0000000000000000000000000000000000000000000000000000000000011000;
    FSM_shift_rows_0_t18 = FSM_shift_rows_0_t17[6'b0 * 1 +: 6 * 1];
    FSM_shift_rows_0_t0[9 * 64 +: 64] = (i_higher_bits >> FSM_shift_rows_0_t18) & 64'b0000000000000000000000000000000000000000000000000000000011111111;
    FSM_shift_rows_0_t0[10 * 64 +: 64] = i_higher_bits & 64'b0000000000000000000000000000000000000000000000000000000011111111;
    FSM_shift_rows_0_t19 = 64'b0000000000000000000000000000000000000000000000000000000000001000;
    FSM_shift_rows_0_t20 = FSM_shift_rows_0_t19[6'b0 * 1 +: 6 * 1];
    FSM_shift_rows_0_t0[11 * 64 +: 64] = (i_higher_bits >> FSM_shift_rows_0_t20) & 64'b0000000000000000000000000000000000000000000000000000000011111111;
    FSM_shift_rows_0_t21 = 64'b0000000000000000000000000000000000000000000000000000000000111000;
    FSM_shift_rows_0_t22 = FSM_shift_rows_0_t21[6'b0 * 1 +: 6 * 1];
    FSM_shift_rows_0_t0[12 * 64 +: 64] = (i_higher_bits >> FSM_shift_rows_0_t22) & 64'b0000000000000000000000000000000000000000000000000000000011111111;
    FSM_shift_rows_0_t23 = 64'b0000000000000000000000000000000000000000000000000000000000100000;
    FSM_shift_rows_0_t24 = FSM_shift_rows_0_t23[6'b0 * 1 +: 6 * 1];
    FSM_shift_rows_0_t0[13 * 64 +: 64] = (i_higher_bits >> FSM_shift_rows_0_t24) & 64'b0000000000000000000000000000000000000000000000000000000011111111;
    FSM_shift_rows_0_t25 = 64'b0000000000000000000000000000000000000000000000000000000000101000;
    FSM_shift_rows_0_t26 = FSM_shift_rows_0_t25[6'b0 * 1 +: 6 * 1];
    FSM_shift_rows_0_t0[14 * 64 +: 64] = (i_higher_bits >> FSM_shift_rows_0_t26) & 64'b0000000000000000000000000000000000000000000000000000000011111111;
    FSM_shift_rows_0_t27 = 64'b0000000000000000000000000000000000000000000000000000000000110000;
    FSM_shift_rows_0_t28 = FSM_shift_rows_0_t27[6'b0 * 1 +: 6 * 1];
    FSM_shift_rows_0_t0[15 * 64 +: 64] = (i_higher_bits >> FSM_shift_rows_0_t28) & 64'b0000000000000000000000000000000000000000000000000000000011111111;
    FSM_shift_rows_0_t29 = 64'b0;
    FSM_shift_rows_0_t30 = FSM_shift_rows_0_t29[6'b0 * 1 +: 4 * 1];
    FSM_shift_rows_0_t31 = FSM_shift_rows_0_t0[FSM_shift_rows_0_t30 * 64 +: 64];
    FSM_shift_rows_0_t32 = 64'b0000000000000000000000000000000000000000000000000000000000111000;
    FSM_shift_rows_0_t33 = FSM_shift_rows_0_t32[6'b0 * 1 +: 6 * 1];
    FSM_shift_rows_0_t34 = 64'b0000000000000000000000000000000000000000000000000000000000000001;
    FSM_shift_rows_0_t35 = FSM_shift_rows_0_t34[6'b0 * 1 +: 4 * 1];
    FSM_shift_rows_0_t36 = FSM_shift_rows_0_t0[FSM_shift_rows_0_t35 * 64 +: 64];
    FSM_shift_rows_0_t37 = 64'b0000000000000000000000000000000000000000000000000000000000110000;
    FSM_shift_rows_0_t38 = FSM_shift_rows_0_t37[6'b0 * 1 +: 6 * 1];
    FSM_shift_rows_0_t39 = 64'b0000000000000000000000000000000000000000000000000000000000000010;
    FSM_shift_rows_0_t40 = FSM_shift_rows_0_t39[6'b0 * 1 +: 4 * 1];
    FSM_shift_rows_0_t41 = FSM_shift_rows_0_t0[FSM_shift_rows_0_t40 * 64 +: 64];
    FSM_shift_rows_0_t42 = 64'b0000000000000000000000000000000000000000000000000000000000101000;
    FSM_shift_rows_0_t43 = FSM_shift_rows_0_t42[6'b0 * 1 +: 6 * 1];
    FSM_shift_rows_0_t44 = 64'b0000000000000000000000000000000000000000000000000000000000000011;
    FSM_shift_rows_0_t45 = FSM_shift_rows_0_t44[6'b0 * 1 +: 4 * 1];
    FSM_shift_rows_0_t46 = FSM_shift_rows_0_t0[FSM_shift_rows_0_t45 * 64 +: 64];
    FSM_shift_rows_0_t47 = 64'b0000000000000000000000000000000000000000000000000000000000100000;
    FSM_shift_rows_0_t48 = FSM_shift_rows_0_t47[6'b0 * 1 +: 6 * 1];
    FSM_shift_rows_0_t49 = 64'b0000000000000000000000000000000000000000000000000000000000000100;
    FSM_shift_rows_0_t50 = FSM_shift_rows_0_t49[6'b0 * 1 +: 4 * 1];
    FSM_shift_rows_0_t51 = FSM_shift_rows_0_t0[FSM_shift_rows_0_t50 * 64 +: 64];
    FSM_shift_rows_0_t52 = 64'b0000000000000000000000000000000000000000000000000000000000011000;
    FSM_shift_rows_0_t53 = FSM_shift_rows_0_t52[6'b0 * 1 +: 6 * 1];
    FSM_shift_rows_0_t54 = 64'b0000000000000000000000000000000000000000000000000000000000000101;
    FSM_shift_rows_0_t55 = FSM_shift_rows_0_t54[6'b0 * 1 +: 4 * 1];
    FSM_shift_rows_0_t56 = FSM_shift_rows_0_t0[FSM_shift_rows_0_t55 * 64 +: 64];
    FSM_shift_rows_0_t57 = 64'b0000000000000000000000000000000000000000000000000000000000010000;
    FSM_shift_rows_0_t58 = FSM_shift_rows_0_t57[6'b0 * 1 +: 6 * 1];
    FSM_shift_rows_0_t59 = 64'b0000000000000000000000000000000000000000000000000000000000000110;
    FSM_shift_rows_0_t60 = FSM_shift_rows_0_t59[6'b0 * 1 +: 4 * 1];
    FSM_shift_rows_0_t61 = FSM_shift_rows_0_t0[FSM_shift_rows_0_t60 * 64 +: 64];
    FSM_shift_rows_0_t62 = 64'b0000000000000000000000000000000000000000000000000000000000001000;
    FSM_shift_rows_0_t63 = FSM_shift_rows_0_t62[6'b0 * 1 +: 6 * 1];
    FSM_shift_rows_0_t64 = 64'b0000000000000000000000000000000000000000000000000000000000000111;
    FSM_shift_rows_0_t65 = FSM_shift_rows_0_t64[6'b0 * 1 +: 4 * 1];
    FSM_shift_rows_0_t66 = FSM_shift_rows_0_t0[FSM_shift_rows_0_t65 * 64 +: 64];
    FSM_shift_rows_0_t67 = 64'b0000000000000000000000000000000000000000000000000000000000001000;
    FSM_shift_rows_0_t68 = FSM_shift_rows_0_t67[6'b0 * 1 +: 4 * 1];
    FSM_shift_rows_0_t69 = FSM_shift_rows_0_t0[FSM_shift_rows_0_t68 * 64 +: 64];
    FSM_shift_rows_0_t70 = 64'b0000000000000000000000000000000000000000000000000000000000111000;
    FSM_shift_rows_0_t71 = FSM_shift_rows_0_t70[6'b0 * 1 +: 6 * 1];
    FSM_shift_rows_0_t72 = 64'b0000000000000000000000000000000000000000000000000000000000001001;
    FSM_shift_rows_0_t73 = FSM_shift_rows_0_t72[6'b0 * 1 +: 4 * 1];
    FSM_shift_rows_0_t74 = FSM_shift_rows_0_t0[FSM_shift_rows_0_t73 * 64 +: 64];
    FSM_shift_rows_0_t75 = 64'b0000000000000000000000000000000000000000000000000000000000110000;
    FSM_shift_rows_0_t76 = FSM_shift_rows_0_t75[6'b0 * 1 +: 6 * 1];
    FSM_shift_rows_0_t77 = 64'b0000000000000000000000000000000000000000000000000000000000001010;
    FSM_shift_rows_0_t78 = FSM_shift_rows_0_t77[6'b0 * 1 +: 4 * 1];
    FSM_shift_rows_0_t79 = FSM_shift_rows_0_t0[FSM_shift_rows_0_t78 * 64 +: 64];
    FSM_shift_rows_0_t80 = 64'b0000000000000000000000000000000000000000000000000000000000101000;
    FSM_shift_rows_0_t81 = FSM_shift_rows_0_t80[6'b0 * 1 +: 6 * 1];
    FSM_shift_rows_0_t82 = 64'b0000000000000000000000000000000000000000000000000000000000001011;
    FSM_shift_rows_0_t83 = FSM_shift_rows_0_t82[6'b0 * 1 +: 4 * 1];
    FSM_shift_rows_0_t84 = FSM_shift_rows_0_t0[FSM_shift_rows_0_t83 * 64 +: 64];
    FSM_shift_rows_0_t85 = 64'b0000000000000000000000000000000000000000000000000000000000100000;
    FSM_shift_rows_0_t86 = FSM_shift_rows_0_t85[6'b0 * 1 +: 6 * 1];
    FSM_shift_rows_0_t87 = 64'b0000000000000000000000000000000000000000000000000000000000001100;
    FSM_shift_rows_0_t88 = FSM_shift_rows_0_t87[6'b0 * 1 +: 4 * 1];
    FSM_shift_rows_0_t89 = FSM_shift_rows_0_t0[FSM_shift_rows_0_t88 * 64 +: 64];
    FSM_shift_rows_0_t90 = 64'b0000000000000000000000000000000000000000000000000000000000011000;
    FSM_shift_rows_0_t91 = FSM_shift_rows_0_t90[6'b0 * 1 +: 6 * 1];
    FSM_shift_rows_0_t92 = 64'b0000000000000000000000000000000000000000000000000000000000001101;
    FSM_shift_rows_0_t93 = FSM_shift_rows_0_t92[6'b0 * 1 +: 4 * 1];
    FSM_shift_rows_0_t94 = FSM_shift_rows_0_t0[FSM_shift_rows_0_t93 * 64 +: 64];
    FSM_shift_rows_0_t95 = 64'b0000000000000000000000000000000000000000000000000000000000010000;
    FSM_shift_rows_0_t96 = FSM_shift_rows_0_t95[6'b0 * 1 +: 6 * 1];
    FSM_shift_rows_0_t97 = 64'b0000000000000000000000000000000000000000000000000000000000001110;
    FSM_shift_rows_0_t98 = FSM_shift_rows_0_t97[6'b0 * 1 +: 4 * 1];
    FSM_shift_rows_0_t99 = FSM_shift_rows_0_t0[FSM_shift_rows_0_t98 * 64 +: 64];
    FSM_shift_rows_0_t100 = 64'b0000000000000000000000000000000000000000000000000000000000001000;
    FSM_shift_rows_0_t101 = FSM_shift_rows_0_t100[6'b0 * 1 +: 6 * 1];
    FSM_shift_rows_0_t102 = 64'b0000000000000000000000000000000000000000000000000000000000001111;
    FSM_shift_rows_0_t103 = FSM_shift_rows_0_t102[6'b0 * 1 +: 4 * 1];
    FSM_shift_rows_0_t104 = FSM_shift_rows_0_t0[FSM_shift_rows_0_t103 * 64 +: 64];
end

always @* begin
    FSM_shift_rows_0_t0[0 * 64 +: 64] = i_lower_bits & 64'b0000000000000000000000000000000000000000000000000000000011111111;
    FSM_shift_rows_0_t1 = 64'b0000000000000000000000000000000000000000000000000000000000001000;
    FSM_shift_rows_0_t2 = FSM_shift_rows_0_t1[6'b0 * 1 +: 6 * 1];
    FSM_shift_rows_0_t0[1 * 64 +: 64] = (i_lower_bits >> FSM_shift_rows_0_t2) & 64'b0000000000000000000000000000000000000000000000000000000011111111;
    FSM_shift_rows_0_t3 = 64'b0000000000000000000000000000000000000000000000000000000000010000;
    FSM_shift_rows_0_t4 = FSM_shift_rows_0_t3[6'b0 * 1 +: 6 * 1];
    FSM_shift_rows_0_t0[2 * 64 +: 64] = (i_lower_bits >> FSM_shift_rows_0_t4) & 64'b0000000000000000000000000000000000000000000000000000000011111111;
    FSM_shift_rows_0_t5 = 64'b0000000000000000000000000000000000000000000000000000000000011000;
    FSM_shift_rows_0_t6 = FSM_shift_rows_0_t5[6'b0 * 1 +: 6 * 1];
    FSM_shift_rows_0_t0[3 * 64 +: 64] = (i_lower_bits >> FSM_shift_rows_0_t6) & 64'b0000000000000000000000000000000000000000000000000000000011111111;
    FSM_shift_rows_0_t7 = 64'b0000000000000000000000000000000000000000000000000000000000101000;
    FSM_shift_rows_0_t8 = FSM_shift_rows_0_t7[6'b0 * 1 +: 6 * 1];
    FSM_shift_rows_0_t0[4 * 64 +: 64] = (i_lower_bits >> FSM_shift_rows_0_t8) & 64'b0000000000000000000000000000000000000000000000000000000011111111;
    FSM_shift_rows_0_t9 = 64'b0000000000000000000000000000000000000000000000000000000000110000;
    FSM_shift_rows_0_t10 = FSM_shift_rows_0_t9[6'b0 * 1 +: 6 * 1];
    FSM_shift_rows_0_t0[5 * 64 +: 64] = (i_lower_bits >> FSM_shift_rows_0_t10) & 64'b0000000000000000000000000000000000000000000000000000000011111111;
    FSM_shift_rows_0_t11 = 64'b0000000000000000000000000000000000000000000000000000000000111000;
    FSM_shift_rows_0_t12 = FSM_shift_rows_0_t11[6'b0 * 1 +: 6 * 1];
    FSM_shift_rows_0_t0[6 * 64 +: 64] = (i_lower_bits >> FSM_shift_rows_0_t12) & 64'b0000000000000000000000000000000000000000000000000000000011111111;
    FSM_shift_rows_0_t13 = 64'b0000000000000000000000000000000000000000000000000000000000100000;
    FSM_shift_rows_0_t14 = FSM_shift_rows_0_t13[6'b0 * 1 +: 6 * 1];
    FSM_shift_rows_0_t0[7 * 64 +: 64] = (i_lower_bits >> FSM_shift_rows_0_t14) & 64'b0000000000000000000000000000000000000000000000000000000011111111;
    FSM_shift_rows_0_t15 = 64'b0000000000000000000000000000000000000000000000000000000000010000;
    FSM_shift_rows_0_t16 = FSM_shift_rows_0_t15[6'b0 * 1 +: 6 * 1];
    FSM_shift_rows_0_t0[8 * 64 +: 64] = (i_higher_bits >> FSM_shift_rows_0_t16) & 64'b0000000000000000000000000000000000000000000000000000000011111111;
    FSM_shift_rows_0_t17 = 64'b0000000000000000000000000000000000000000000000000000000000011000;
    FSM_shift_rows_0_t18 = FSM_shift_rows_0_t17[6'b0 * 1 +: 6 * 1];
    FSM_shift_rows_0_t0[9 * 64 +: 64] = (i_higher_bits >> FSM_shift_rows_0_t18) & 64'b0000000000000000000000000000000000000000000000000000000011111111;
    FSM_shift_rows_0_t0[10 * 64 +: 64] = i_higher_bits & 64'b0000000000000000000000000000000000000000000000000000000011111111;
    FSM_shift_rows_0_t19 = 64'b0000000000000000000000000000000000000000000000000000000000001000;
    FSM_shift_rows_0_t20 = FSM_shift_rows_0_t19[6'b0 * 1 +: 6 * 1];
    FSM_shift_rows_0_t0[11 * 64 +: 64] = (i_higher_bits >> FSM_shift_rows_0_t20) & 64'b0000000000000000000000000000000000000000000000000000000011111111;
    FSM_shift_rows_0_t21 = 64'b0000000000000000000000000000000000000000000000000000000000111000;
    FSM_shift_rows_0_t22 = FSM_shift_rows_0_t21[6'b0 * 1 +: 6 * 1];
    FSM_shift_rows_0_t0[12 * 64 +: 64] = (i_higher_bits >> FSM_shift_rows_0_t22) & 64'b0000000000000000000000000000000000000000000000000000000011111111;
    FSM_shift_rows_0_t23 = 64'b0000000000000000000000000000000000000000000000000000000000100000;
    FSM_shift_rows_0_t24 = FSM_shift_rows_0_t23[6'b0 * 1 +: 6 * 1];
    FSM_shift_rows_0_t0[13 * 64 +: 64] = (i_higher_bits >> FSM_shift_rows_0_t24) & 64'b0000000000000000000000000000000000000000000000000000000011111111;
    FSM_shift_rows_0_t25 = 64'b0000000000000000000000000000000000000000000000000000000000101000;
    FSM_shift_rows_0_t26 = FSM_shift_rows_0_t25[6'b0 * 1 +: 6 * 1];
    FSM_shift_rows_0_t0[14 * 64 +: 64] = (i_higher_bits >> FSM_shift_rows_0_t26) & 64'b0000000000000000000000000000000000000000000000000000000011111111;
    FSM_shift_rows_0_t27 = 64'b0000000000000000000000000000000000000000000000000000000000110000;
    FSM_shift_rows_0_t28 = FSM_shift_rows_0_t27[6'b0 * 1 +: 6 * 1];
    FSM_shift_rows_0_t0[15 * 64 +: 64] = (i_higher_bits >> FSM_shift_rows_0_t28) & 64'b0000000000000000000000000000000000000000000000000000000011111111;
    FSM_shift_rows_0_t29 = 64'b0;
    FSM_shift_rows_0_t30 = FSM_shift_rows_0_t29[6'b0 * 1 +: 4 * 1];
    FSM_shift_rows_0_t31 = FSM_shift_rows_0_t0[FSM_shift_rows_0_t30 * 64 +: 64];
    FSM_shift_rows_0_t32 = 64'b0000000000000000000000000000000000000000000000000000000000111000;
    FSM_shift_rows_0_t33 = FSM_shift_rows_0_t32[6'b0 * 1 +: 6 * 1];
    FSM_shift_rows_0_t34 = 64'b0000000000000000000000000000000000000000000000000000000000000001;
    FSM_shift_rows_0_t35 = FSM_shift_rows_0_t34[6'b0 * 1 +: 4 * 1];
    FSM_shift_rows_0_t36 = FSM_shift_rows_0_t0[FSM_shift_rows_0_t35 * 64 +: 64];
    FSM_shift_rows_0_t37 = 64'b0000000000000000000000000000000000000000000000000000000000110000;
    FSM_shift_rows_0_t38 = FSM_shift_rows_0_t37[6'b0 * 1 +: 6 * 1];
    FSM_shift_rows_0_t39 = 64'b0000000000000000000000000000000000000000000000000000000000000010;
    FSM_shift_rows_0_t40 = FSM_shift_rows_0_t39[6'b0 * 1 +: 4 * 1];
    FSM_shift_rows_0_t41 = FSM_shift_rows_0_t0[FSM_shift_rows_0_t40 * 64 +: 64];
    FSM_shift_rows_0_t42 = 64'b0000000000000000000000000000000000000000000000000000000000101000;
    FSM_shift_rows_0_t43 = FSM_shift_rows_0_t42[6'b0 * 1 +: 6 * 1];
    FSM_shift_rows_0_t44 = 64'b0000000000000000000000000000000000000000000000000000000000000011;
    FSM_shift_rows_0_t45 = FSM_shift_rows_0_t44[6'b0 * 1 +: 4 * 1];
    FSM_shift_rows_0_t46 = FSM_shift_rows_0_t0[FSM_shift_rows_0_t45 * 64 +: 64];
    FSM_shift_rows_0_t47 = 64'b0000000000000000000000000000000000000000000000000000000000100000;
    FSM_shift_rows_0_t48 = FSM_shift_rows_0_t47[6'b0 * 1 +: 6 * 1];
    FSM_shift_rows_0_t49 = 64'b0000000000000000000000000000000000000000000000000000000000000100;
    FSM_shift_rows_0_t50 = FSM_shift_rows_0_t49[6'b0 * 1 +: 4 * 1];
    FSM_shift_rows_0_t51 = FSM_shift_rows_0_t0[FSM_shift_rows_0_t50 * 64 +: 64];
    FSM_shift_rows_0_t52 = 64'b0000000000000000000000000000000000000000000000000000000000011000;
    FSM_shift_rows_0_t53 = FSM_shift_rows_0_t52[6'b0 * 1 +: 6 * 1];
    FSM_shift_rows_0_t54 = 64'b0000000000000000000000000000000000000000000000000000000000000101;
    FSM_shift_rows_0_t55 = FSM_shift_rows_0_t54[6'b0 * 1 +: 4 * 1];
    FSM_shift_rows_0_t56 = FSM_shift_rows_0_t0[FSM_shift_rows_0_t55 * 64 +: 64];
    FSM_shift_rows_0_t57 = 64'b0000000000000000000000000000000000000000000000000000000000010000;
    FSM_shift_rows_0_t58 = FSM_shift_rows_0_t57[6'b0 * 1 +: 6 * 1];
    FSM_shift_rows_0_t59 = 64'b0000000000000000000000000000000000000000000000000000000000000110;
    FSM_shift_rows_0_t60 = FSM_shift_rows_0_t59[6'b0 * 1 +: 4 * 1];
    FSM_shift_rows_0_t61 = FSM_shift_rows_0_t0[FSM_shift_rows_0_t60 * 64 +: 64];
    FSM_shift_rows_0_t62 = 64'b0000000000000000000000000000000000000000000000000000000000001000;
    FSM_shift_rows_0_t63 = FSM_shift_rows_0_t62[6'b0 * 1 +: 6 * 1];
    FSM_shift_rows_0_t64 = 64'b0000000000000000000000000000000000000000000000000000000000000111;
    FSM_shift_rows_0_t65 = FSM_shift_rows_0_t64[6'b0 * 1 +: 4 * 1];
    FSM_shift_rows_0_t66 = FSM_shift_rows_0_t0[FSM_shift_rows_0_t65 * 64 +: 64];
    FSM_shift_rows_0_t67 = 64'b0000000000000000000000000000000000000000000000000000000000001000;
    FSM_shift_rows_0_t68 = FSM_shift_rows_0_t67[6'b0 * 1 +: 4 * 1];
    FSM_shift_rows_0_t69 = FSM_shift_rows_0_t0[FSM_shift_rows_0_t68 * 64 +: 64];
    FSM_shift_rows_0_t70 = 64'b0000000000000000000000000000000000000000000000000000000000111000;
    FSM_shift_rows_0_t71 = FSM_shift_rows_0_t70[6'b0 * 1 +: 6 * 1];
    FSM_shift_rows_0_t72 = 64'b0000000000000000000000000000000000000000000000000000000000001001;
    FSM_shift_rows_0_t73 = FSM_shift_rows_0_t72[6'b0 * 1 +: 4 * 1];
    FSM_shift_rows_0_t74 = FSM_shift_rows_0_t0[FSM_shift_rows_0_t73 * 64 +: 64];
    FSM_shift_rows_0_t75 = 64'b0000000000000000000000000000000000000000000000000000000000110000;
    FSM_shift_rows_0_t76 = FSM_shift_rows_0_t75[6'b0 * 1 +: 6 * 1];
    FSM_shift_rows_0_t77 = 64'b0000000000000000000000000000000000000000000000000000000000001010;
    FSM_shift_rows_0_t78 = FSM_shift_rows_0_t77[6'b0 * 1 +: 4 * 1];
    FSM_shift_rows_0_t79 = FSM_shift_rows_0_t0[FSM_shift_rows_0_t78 * 64 +: 64];
    FSM_shift_rows_0_t80 = 64'b0000000000000000000000000000000000000000000000000000000000101000;
    FSM_shift_rows_0_t81 = FSM_shift_rows_0_t80[6'b0 * 1 +: 6 * 1];
    FSM_shift_rows_0_t82 = 64'b0000000000000000000000000000000000000000000000000000000000001011;
    FSM_shift_rows_0_t83 = FSM_shift_rows_0_t82[6'b0 * 1 +: 4 * 1];
    FSM_shift_rows_0_t84 = FSM_shift_rows_0_t0[FSM_shift_rows_0_t83 * 64 +: 64];
    FSM_shift_rows_0_t85 = 64'b0000000000000000000000000000000000000000000000000000000000100000;
    FSM_shift_rows_0_t86 = FSM_shift_rows_0_t85[6'b0 * 1 +: 6 * 1];
    FSM_shift_rows_0_t87 = 64'b0000000000000000000000000000000000000000000000000000000000001100;
    FSM_shift_rows_0_t88 = FSM_shift_rows_0_t87[6'b0 * 1 +: 4 * 1];
    FSM_shift_rows_0_t89 = FSM_shift_rows_0_t0[FSM_shift_rows_0_t88 * 64 +: 64];
    FSM_shift_rows_0_t90 = 64'b0000000000000000000000000000000000000000000000000000000000011000;
    FSM_shift_rows_0_t91 = FSM_shift_rows_0_t90[6'b0 * 1 +: 6 * 1];
    FSM_shift_rows_0_t92 = 64'b0000000000000000000000000000000000000000000000000000000000001101;
    FSM_shift_rows_0_t93 = FSM_shift_rows_0_t92[6'b0 * 1 +: 4 * 1];
    FSM_shift_rows_0_t94 = FSM_shift_rows_0_t0[FSM_shift_rows_0_t93 * 64 +: 64];
    FSM_shift_rows_0_t95 = 64'b0000000000000000000000000000000000000000000000000000000000010000;
    FSM_shift_rows_0_t96 = FSM_shift_rows_0_t95[6'b0 * 1 +: 6 * 1];
    FSM_shift_rows_0_t97 = 64'b0000000000000000000000000000000000000000000000000000000000001110;
    FSM_shift_rows_0_t98 = FSM_shift_rows_0_t97[6'b0 * 1 +: 4 * 1];
    FSM_shift_rows_0_t99 = FSM_shift_rows_0_t0[FSM_shift_rows_0_t98 * 64 +: 64];
    FSM_shift_rows_0_t100 = 64'b0000000000000000000000000000000000000000000000000000000000001000;
    FSM_shift_rows_0_t101 = FSM_shift_rows_0_t100[6'b0 * 1 +: 6 * 1];
    FSM_shift_rows_0_t102 = 64'b0000000000000000000000000000000000000000000000000000000000001111;
    FSM_shift_rows_0_t103 = FSM_shift_rows_0_t102[6'b0 * 1 +: 4 * 1];
    FSM_shift_rows_0_t104 = FSM_shift_rows_0_t0[FSM_shift_rows_0_t103 * 64 +: 64];
end

assign FSM_shift_rows_0_in_ready = 1'b1;

always @(posedge clk) begin
    FSM_shift_rows_0_st_dummy_reg <= FSM_shift_rows_0_st_dummy_reg;
    if (rst) begin
        FSM_shift_rows_0_st_dummy_reg <= 64'b0;
    end
end
/* End submodules of shift_rows */
/* End module shift_rows */
endgenerate
endmodule
