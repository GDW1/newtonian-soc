`timescale 1ns / 1ps

module dct_8x8_stage_7_inner
(
    input wire clk,
    input wire rst,
    input wire [2048-1:0] i_data_in,
    input wire i_valid,
    output wire i_ready,
    output wire [2048-1:0] o_data_out,
    output wire o_valid,
    input wire o_ready
);

generate
/*
    Begin module dct_8x8_stage_7
*/
/*
    Wires declared by dct_8x8_stage_7
*/
wire FSM_dct_8x8_stage_7_0_in_ready;
wire FSM_dct_8x8_stage_7_0_out_valid;
/* End wires declared by dct_8x8_stage_7 */

/*
    Submodules of dct_8x8_stage_7
*/
reg [32-1:0] FSM_dct_8x8_stage_7_0_st_dummy_reg = 32'b0;

reg [32-1:0] FSM_dct_8x8_stage_7_0_t0;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t1;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t2;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t3;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t4;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t5;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t6;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t7;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t8;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t9;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t10;
reg [2048-1:0] FSM_dct_8x8_stage_7_0_t11;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t12;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t13;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t14;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t15;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t16;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t17;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t18;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t19;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t20;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t21;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t22;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t23;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t24;
reg [2048-1:0] FSM_dct_8x8_stage_7_0_t25;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t26;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t27;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t28;
reg [2048-1:0] FSM_dct_8x8_stage_7_0_t29;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t30;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t31;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t32;
reg [2048-1:0] FSM_dct_8x8_stage_7_0_t33;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t34;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t35;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t36;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t37;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t38;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t39;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t40;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t41;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t42;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t43;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t44;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t45;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t46;
reg [2048-1:0] FSM_dct_8x8_stage_7_0_t47;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t48;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t49;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t50;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t51;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t52;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t53;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t54;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t55;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t56;
reg [2048-1:0] FSM_dct_8x8_stage_7_0_t57;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t58;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t59;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t60;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t61;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t62;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t63;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t64;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t65;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t66;
reg [2048-1:0] FSM_dct_8x8_stage_7_0_t67;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t68;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t69;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t70;
reg [2048-1:0] FSM_dct_8x8_stage_7_0_t71;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t72;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t73;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t74;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t75;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t76;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t77;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t78;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t79;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t80;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t81;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t82;
reg [2048-1:0] FSM_dct_8x8_stage_7_0_t83;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t84;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t85;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t86;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t87;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t88;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t89;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t90;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t91;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t92;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t93;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t94;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t95;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t96;
reg [2048-1:0] FSM_dct_8x8_stage_7_0_t97;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t98;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t99;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t100;
reg [2048-1:0] FSM_dct_8x8_stage_7_0_t101;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t102;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t103;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t104;
reg [2048-1:0] FSM_dct_8x8_stage_7_0_t105;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t106;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t107;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t108;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t109;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t110;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t111;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t112;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t113;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t114;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t115;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t116;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t117;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t118;
reg [2048-1:0] FSM_dct_8x8_stage_7_0_t119;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t120;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t121;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t122;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t123;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t124;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t125;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t126;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t127;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t128;
reg [2048-1:0] FSM_dct_8x8_stage_7_0_t129;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t130;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t131;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t132;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t133;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t134;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t135;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t136;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t137;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t138;
reg [2048-1:0] FSM_dct_8x8_stage_7_0_t139;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t140;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t141;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t142;
reg [2048-1:0] FSM_dct_8x8_stage_7_0_t143;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t144;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t145;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t146;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t147;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t148;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t149;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t150;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t151;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t152;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t153;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t154;
reg [2048-1:0] FSM_dct_8x8_stage_7_0_t155;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t156;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t157;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t158;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t159;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t160;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t161;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t162;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t163;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t164;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t165;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t166;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t167;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t168;
reg [2048-1:0] FSM_dct_8x8_stage_7_0_t169;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t170;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t171;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t172;
reg [2048-1:0] FSM_dct_8x8_stage_7_0_t173;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t174;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t175;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t176;
reg [2048-1:0] FSM_dct_8x8_stage_7_0_t177;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t178;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t179;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t180;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t181;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t182;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t183;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t184;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t185;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t186;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t187;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t188;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t189;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t190;
reg [2048-1:0] FSM_dct_8x8_stage_7_0_t191;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t192;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t193;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t194;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t195;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t196;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t197;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t198;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t199;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t200;
reg [2048-1:0] FSM_dct_8x8_stage_7_0_t201;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t202;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t203;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t204;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t205;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t206;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t207;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t208;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t209;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t210;
reg [2048-1:0] FSM_dct_8x8_stage_7_0_t211;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t212;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t213;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t214;
reg [2048-1:0] FSM_dct_8x8_stage_7_0_t215;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t216;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t217;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t218;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t219;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t220;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t221;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t222;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t223;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t224;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t225;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t226;
reg [2048-1:0] FSM_dct_8x8_stage_7_0_t227;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t228;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t229;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t230;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t231;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t232;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t233;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t234;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t235;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t236;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t237;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t238;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t239;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t240;
reg [2048-1:0] FSM_dct_8x8_stage_7_0_t241;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t242;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t243;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t244;
reg [2048-1:0] FSM_dct_8x8_stage_7_0_t245;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t246;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t247;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t248;
reg [2048-1:0] FSM_dct_8x8_stage_7_0_t249;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t250;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t251;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t252;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t253;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t254;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t255;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t256;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t257;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t258;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t259;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t260;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t261;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t262;
reg [2048-1:0] FSM_dct_8x8_stage_7_0_t263;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t264;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t265;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t266;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t267;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t268;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t269;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t270;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t271;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t272;
reg [2048-1:0] FSM_dct_8x8_stage_7_0_t273;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t274;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t275;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t276;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t277;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t278;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t279;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t280;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t281;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t282;
reg [2048-1:0] FSM_dct_8x8_stage_7_0_t283;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t284;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t285;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t286;
reg [2048-1:0] FSM_dct_8x8_stage_7_0_t287;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t288;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t289;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t290;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t291;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t292;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t293;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t294;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t295;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t296;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t297;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t298;
reg [2048-1:0] FSM_dct_8x8_stage_7_0_t299;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t300;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t301;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t302;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t303;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t304;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t305;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t306;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t307;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t308;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t309;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t310;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t311;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t312;
reg [2048-1:0] FSM_dct_8x8_stage_7_0_t313;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t314;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t315;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t316;
reg [2048-1:0] FSM_dct_8x8_stage_7_0_t317;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t318;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t319;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t320;
reg [2048-1:0] FSM_dct_8x8_stage_7_0_t321;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t322;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t323;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t324;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t325;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t326;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t327;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t328;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t329;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t330;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t331;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t332;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t333;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t334;
reg [2048-1:0] FSM_dct_8x8_stage_7_0_t335;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t336;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t337;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t338;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t339;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t340;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t341;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t342;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t343;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t344;
reg [2048-1:0] FSM_dct_8x8_stage_7_0_t345;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t346;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t347;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t348;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t349;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t350;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t351;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t352;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t353;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t354;
reg [2048-1:0] FSM_dct_8x8_stage_7_0_t355;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t356;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t357;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t358;
reg [2048-1:0] FSM_dct_8x8_stage_7_0_t359;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t360;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t361;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t362;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t363;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t364;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t365;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t366;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t367;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t368;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t369;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t370;
reg [2048-1:0] FSM_dct_8x8_stage_7_0_t371;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t372;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t373;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t374;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t375;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t376;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t377;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t378;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t379;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t380;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t381;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t382;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t383;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t384;
reg [2048-1:0] FSM_dct_8x8_stage_7_0_t385;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t386;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t387;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t388;
reg [2048-1:0] FSM_dct_8x8_stage_7_0_t389;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t390;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t391;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t392;
reg [2048-1:0] FSM_dct_8x8_stage_7_0_t393;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t394;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t395;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t396;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t397;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t398;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t399;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t400;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t401;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t402;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t403;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t404;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t405;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t406;
reg [2048-1:0] FSM_dct_8x8_stage_7_0_t407;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t408;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t409;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t410;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t411;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t412;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t413;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t414;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t415;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t416;
reg [2048-1:0] FSM_dct_8x8_stage_7_0_t417;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t418;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t419;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t420;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t421;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t422;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t423;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t424;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t425;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t426;
reg [2048-1:0] FSM_dct_8x8_stage_7_0_t427;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t428;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t429;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t430;
reg [2048-1:0] FSM_dct_8x8_stage_7_0_t431;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t432;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t433;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t434;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t435;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t436;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t437;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t438;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t439;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t440;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t441;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t442;
reg [2048-1:0] FSM_dct_8x8_stage_7_0_t443;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t444;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t445;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t446;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t447;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t448;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t449;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t450;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t451;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t452;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t453;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t454;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t455;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t456;
reg [2048-1:0] FSM_dct_8x8_stage_7_0_t457;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t458;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t459;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t460;
reg [2048-1:0] FSM_dct_8x8_stage_7_0_t461;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t462;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t463;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t464;
reg [2048-1:0] FSM_dct_8x8_stage_7_0_t465;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t466;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t467;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t468;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t469;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t470;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t471;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t472;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t473;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t474;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t475;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t476;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t477;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t478;
reg [2048-1:0] FSM_dct_8x8_stage_7_0_t479;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t480;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t481;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t482;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t483;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t484;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t485;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t486;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t487;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t488;
reg [2048-1:0] FSM_dct_8x8_stage_7_0_t489;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t490;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t491;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t492;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t493;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t494;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t495;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t496;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t497;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t498;
reg [2048-1:0] FSM_dct_8x8_stage_7_0_t499;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t500;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t501;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t502;
reg [2048-1:0] FSM_dct_8x8_stage_7_0_t503;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t504;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t505;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t506;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t507;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t508;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t509;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t510;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t511;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t512;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t513;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t514;
reg [2048-1:0] FSM_dct_8x8_stage_7_0_t515;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t516;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t517;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t518;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t519;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t520;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t521;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t522;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t523;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t524;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t525;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t526;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t527;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t528;
reg [2048-1:0] FSM_dct_8x8_stage_7_0_t529;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t530;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t531;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t532;
reg [2048-1:0] FSM_dct_8x8_stage_7_0_t533;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t534;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t535;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t536;
reg [2048-1:0] FSM_dct_8x8_stage_7_0_t537;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t538;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t539;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t540;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t541;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t542;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t543;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t544;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t545;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t546;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t547;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t548;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t549;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t550;
reg [2048-1:0] FSM_dct_8x8_stage_7_0_t551;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t552;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t553;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t554;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t555;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t556;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t557;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t558;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t559;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t560;
reg [2048-1:0] FSM_dct_8x8_stage_7_0_t561;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t562;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t563;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t564;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t565;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t566;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t567;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t568;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t569;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t570;
reg [2048-1:0] FSM_dct_8x8_stage_7_0_t571;
reg [33-1:0] FSM_dct_8x8_stage_7_0_t572;
reg [32-1:0] FSM_dct_8x8_stage_7_0_t573;
reg [6-1:0] FSM_dct_8x8_stage_7_0_t574;
reg [2048-1:0] FSM_dct_8x8_stage_7_0_t575;

/*
    Wiring by dct_8x8_stage_7
*/
assign i_ready = FSM_dct_8x8_stage_7_0_in_ready;
assign o_data_out = FSM_dct_8x8_stage_7_0_t575;
assign o_valid = FSM_dct_8x8_stage_7_0_out_valid;
/* End wiring by dct_8x8_stage_7 */

assign FSM_dct_8x8_stage_7_0_out_valid = 1'b1;

initial begin
    FSM_dct_8x8_stage_7_0_t0 = 32'b0;
    FSM_dct_8x8_stage_7_0_t1 = FSM_dct_8x8_stage_7_0_t0[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t2 = 32'b0;
    FSM_dct_8x8_stage_7_0_t3 = FSM_dct_8x8_stage_7_0_t2[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t4 = i_data_in[FSM_dct_8x8_stage_7_0_t3 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t5 = 32'b00000000000000000000000000011000 + 32'b0;
    FSM_dct_8x8_stage_7_0_t6 = FSM_dct_8x8_stage_7_0_t5[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t7 = FSM_dct_8x8_stage_7_0_t6[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t8 = i_data_in[FSM_dct_8x8_stage_7_0_t7 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t9 = FSM_dct_8x8_stage_7_0_t4 + FSM_dct_8x8_stage_7_0_t8;
    FSM_dct_8x8_stage_7_0_t10 = FSM_dct_8x8_stage_7_0_t9[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t11 = 2048'b0;
    FSM_dct_8x8_stage_7_0_t11[FSM_dct_8x8_stage_7_0_t1 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t10;
    FSM_dct_8x8_stage_7_0_t12 = 32'b00000000000000000000000000001000 + 32'b0;
    FSM_dct_8x8_stage_7_0_t13 = FSM_dct_8x8_stage_7_0_t12[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t14 = FSM_dct_8x8_stage_7_0_t13[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t15 = 32'b00000000000000000000000000001000 + 32'b0;
    FSM_dct_8x8_stage_7_0_t16 = FSM_dct_8x8_stage_7_0_t15[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t17 = FSM_dct_8x8_stage_7_0_t16[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t18 = i_data_in[FSM_dct_8x8_stage_7_0_t17 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t19 = 32'b00000000000000000000000000010000 + 32'b0;
    FSM_dct_8x8_stage_7_0_t20 = FSM_dct_8x8_stage_7_0_t19[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t21 = FSM_dct_8x8_stage_7_0_t20[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t22 = i_data_in[FSM_dct_8x8_stage_7_0_t21 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t23 = FSM_dct_8x8_stage_7_0_t18 + FSM_dct_8x8_stage_7_0_t22;
    FSM_dct_8x8_stage_7_0_t24 = FSM_dct_8x8_stage_7_0_t23[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t25 = FSM_dct_8x8_stage_7_0_t11;
    FSM_dct_8x8_stage_7_0_t25[FSM_dct_8x8_stage_7_0_t14 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t24;
    FSM_dct_8x8_stage_7_0_t26 = 32'b00000000000000000000000000010000 + 32'b0;
    FSM_dct_8x8_stage_7_0_t27 = FSM_dct_8x8_stage_7_0_t26[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t28 = FSM_dct_8x8_stage_7_0_t27[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t29 = FSM_dct_8x8_stage_7_0_t25;
    FSM_dct_8x8_stage_7_0_t29[FSM_dct_8x8_stage_7_0_t28 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t18 - FSM_dct_8x8_stage_7_0_t22;
    FSM_dct_8x8_stage_7_0_t30 = 32'b00000000000000000000000000011000 + 32'b0;
    FSM_dct_8x8_stage_7_0_t31 = FSM_dct_8x8_stage_7_0_t30[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t32 = FSM_dct_8x8_stage_7_0_t31[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t33 = FSM_dct_8x8_stage_7_0_t29;
    FSM_dct_8x8_stage_7_0_t33[FSM_dct_8x8_stage_7_0_t32 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t4 - FSM_dct_8x8_stage_7_0_t8;
    FSM_dct_8x8_stage_7_0_t34 = 32'b00000000000000000000000000100000 + 32'b0;
    FSM_dct_8x8_stage_7_0_t35 = FSM_dct_8x8_stage_7_0_t34[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t36 = FSM_dct_8x8_stage_7_0_t35[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t37 = 32'b00000000000000000000000000100000 + 32'b0;
    FSM_dct_8x8_stage_7_0_t38 = FSM_dct_8x8_stage_7_0_t37[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t39 = FSM_dct_8x8_stage_7_0_t38[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t40 = i_data_in[FSM_dct_8x8_stage_7_0_t39 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t41 = 32'b00000000000000000000000000101000 + 32'b0;
    FSM_dct_8x8_stage_7_0_t42 = FSM_dct_8x8_stage_7_0_t41[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t43 = FSM_dct_8x8_stage_7_0_t42[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t44 = i_data_in[FSM_dct_8x8_stage_7_0_t43 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t45 = FSM_dct_8x8_stage_7_0_t40 + FSM_dct_8x8_stage_7_0_t44;
    FSM_dct_8x8_stage_7_0_t46 = FSM_dct_8x8_stage_7_0_t45[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t47 = FSM_dct_8x8_stage_7_0_t33;
    FSM_dct_8x8_stage_7_0_t47[FSM_dct_8x8_stage_7_0_t36 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t46;
    FSM_dct_8x8_stage_7_0_t48 = 32'b00000000000000000000000000101000 + 32'b0;
    FSM_dct_8x8_stage_7_0_t49 = FSM_dct_8x8_stage_7_0_t48[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t50 = FSM_dct_8x8_stage_7_0_t49[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t51 = 32'b00000000000000000000000000110000 + 32'b0;
    FSM_dct_8x8_stage_7_0_t52 = FSM_dct_8x8_stage_7_0_t51[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t53 = FSM_dct_8x8_stage_7_0_t52[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t54 = i_data_in[FSM_dct_8x8_stage_7_0_t53 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t55 = FSM_dct_8x8_stage_7_0_t44 + FSM_dct_8x8_stage_7_0_t54;
    FSM_dct_8x8_stage_7_0_t56 = FSM_dct_8x8_stage_7_0_t55[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t57 = FSM_dct_8x8_stage_7_0_t47;
    FSM_dct_8x8_stage_7_0_t57[FSM_dct_8x8_stage_7_0_t50 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t56;
    FSM_dct_8x8_stage_7_0_t58 = 32'b00000000000000000000000000110000 + 32'b0;
    FSM_dct_8x8_stage_7_0_t59 = FSM_dct_8x8_stage_7_0_t58[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t60 = FSM_dct_8x8_stage_7_0_t59[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t61 = 32'b00000000000000000000000000111000 + 32'b0;
    FSM_dct_8x8_stage_7_0_t62 = FSM_dct_8x8_stage_7_0_t61[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t63 = FSM_dct_8x8_stage_7_0_t62[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t64 = i_data_in[FSM_dct_8x8_stage_7_0_t63 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t65 = FSM_dct_8x8_stage_7_0_t54 + FSM_dct_8x8_stage_7_0_t64;
    FSM_dct_8x8_stage_7_0_t66 = FSM_dct_8x8_stage_7_0_t65[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t67 = FSM_dct_8x8_stage_7_0_t57;
    FSM_dct_8x8_stage_7_0_t67[FSM_dct_8x8_stage_7_0_t60 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t66;
    FSM_dct_8x8_stage_7_0_t68 = 32'b00000000000000000000000000111000 + 32'b0;
    FSM_dct_8x8_stage_7_0_t69 = FSM_dct_8x8_stage_7_0_t68[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t70 = FSM_dct_8x8_stage_7_0_t69[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t71 = FSM_dct_8x8_stage_7_0_t67;
    FSM_dct_8x8_stage_7_0_t71[FSM_dct_8x8_stage_7_0_t70 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t64;
    FSM_dct_8x8_stage_7_0_t72 = 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_7_0_t73 = FSM_dct_8x8_stage_7_0_t72[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t74 = 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_7_0_t75 = FSM_dct_8x8_stage_7_0_t74[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t76 = i_data_in[FSM_dct_8x8_stage_7_0_t75 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t77 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_7_0_t78 = FSM_dct_8x8_stage_7_0_t77[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t79 = FSM_dct_8x8_stage_7_0_t78[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t80 = i_data_in[FSM_dct_8x8_stage_7_0_t79 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t81 = FSM_dct_8x8_stage_7_0_t76 + FSM_dct_8x8_stage_7_0_t80;
    FSM_dct_8x8_stage_7_0_t82 = FSM_dct_8x8_stage_7_0_t81[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t83 = FSM_dct_8x8_stage_7_0_t71;
    FSM_dct_8x8_stage_7_0_t83[FSM_dct_8x8_stage_7_0_t73 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t82;
    FSM_dct_8x8_stage_7_0_t84 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_7_0_t85 = FSM_dct_8x8_stage_7_0_t84[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t86 = FSM_dct_8x8_stage_7_0_t85[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t87 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_7_0_t88 = FSM_dct_8x8_stage_7_0_t87[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t89 = FSM_dct_8x8_stage_7_0_t88[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t90 = i_data_in[FSM_dct_8x8_stage_7_0_t89 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t91 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_7_0_t92 = FSM_dct_8x8_stage_7_0_t91[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t93 = FSM_dct_8x8_stage_7_0_t92[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t94 = i_data_in[FSM_dct_8x8_stage_7_0_t93 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t95 = FSM_dct_8x8_stage_7_0_t90 + FSM_dct_8x8_stage_7_0_t94;
    FSM_dct_8x8_stage_7_0_t96 = FSM_dct_8x8_stage_7_0_t95[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t97 = FSM_dct_8x8_stage_7_0_t83;
    FSM_dct_8x8_stage_7_0_t97[FSM_dct_8x8_stage_7_0_t86 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t96;
    FSM_dct_8x8_stage_7_0_t98 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_7_0_t99 = FSM_dct_8x8_stage_7_0_t98[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t100 = FSM_dct_8x8_stage_7_0_t99[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t101 = FSM_dct_8x8_stage_7_0_t97;
    FSM_dct_8x8_stage_7_0_t101[FSM_dct_8x8_stage_7_0_t100 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t90 - FSM_dct_8x8_stage_7_0_t94;
    FSM_dct_8x8_stage_7_0_t102 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_7_0_t103 = FSM_dct_8x8_stage_7_0_t102[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t104 = FSM_dct_8x8_stage_7_0_t103[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t105 = FSM_dct_8x8_stage_7_0_t101;
    FSM_dct_8x8_stage_7_0_t105[FSM_dct_8x8_stage_7_0_t104 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t76 - FSM_dct_8x8_stage_7_0_t80;
    FSM_dct_8x8_stage_7_0_t106 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_7_0_t107 = FSM_dct_8x8_stage_7_0_t106[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t108 = FSM_dct_8x8_stage_7_0_t107[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t109 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_7_0_t110 = FSM_dct_8x8_stage_7_0_t109[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t111 = FSM_dct_8x8_stage_7_0_t110[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t112 = i_data_in[FSM_dct_8x8_stage_7_0_t111 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t113 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_7_0_t114 = FSM_dct_8x8_stage_7_0_t113[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t115 = FSM_dct_8x8_stage_7_0_t114[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t116 = i_data_in[FSM_dct_8x8_stage_7_0_t115 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t117 = FSM_dct_8x8_stage_7_0_t112 + FSM_dct_8x8_stage_7_0_t116;
    FSM_dct_8x8_stage_7_0_t118 = FSM_dct_8x8_stage_7_0_t117[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t119 = FSM_dct_8x8_stage_7_0_t105;
    FSM_dct_8x8_stage_7_0_t119[FSM_dct_8x8_stage_7_0_t108 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t118;
    FSM_dct_8x8_stage_7_0_t120 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_7_0_t121 = FSM_dct_8x8_stage_7_0_t120[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t122 = FSM_dct_8x8_stage_7_0_t121[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t123 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_7_0_t124 = FSM_dct_8x8_stage_7_0_t123[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t125 = FSM_dct_8x8_stage_7_0_t124[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t126 = i_data_in[FSM_dct_8x8_stage_7_0_t125 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t127 = FSM_dct_8x8_stage_7_0_t116 + FSM_dct_8x8_stage_7_0_t126;
    FSM_dct_8x8_stage_7_0_t128 = FSM_dct_8x8_stage_7_0_t127[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t129 = FSM_dct_8x8_stage_7_0_t119;
    FSM_dct_8x8_stage_7_0_t129[FSM_dct_8x8_stage_7_0_t122 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t128;
    FSM_dct_8x8_stage_7_0_t130 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_7_0_t131 = FSM_dct_8x8_stage_7_0_t130[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t132 = FSM_dct_8x8_stage_7_0_t131[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t133 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_7_0_t134 = FSM_dct_8x8_stage_7_0_t133[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t135 = FSM_dct_8x8_stage_7_0_t134[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t136 = i_data_in[FSM_dct_8x8_stage_7_0_t135 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t137 = FSM_dct_8x8_stage_7_0_t126 + FSM_dct_8x8_stage_7_0_t136;
    FSM_dct_8x8_stage_7_0_t138 = FSM_dct_8x8_stage_7_0_t137[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t139 = FSM_dct_8x8_stage_7_0_t129;
    FSM_dct_8x8_stage_7_0_t139[FSM_dct_8x8_stage_7_0_t132 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t138;
    FSM_dct_8x8_stage_7_0_t140 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_7_0_t141 = FSM_dct_8x8_stage_7_0_t140[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t142 = FSM_dct_8x8_stage_7_0_t141[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t143 = FSM_dct_8x8_stage_7_0_t139;
    FSM_dct_8x8_stage_7_0_t143[FSM_dct_8x8_stage_7_0_t142 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t136;
    FSM_dct_8x8_stage_7_0_t144 = 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_7_0_t145 = FSM_dct_8x8_stage_7_0_t144[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t146 = 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_7_0_t147 = FSM_dct_8x8_stage_7_0_t146[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t148 = i_data_in[FSM_dct_8x8_stage_7_0_t147 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t149 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_7_0_t150 = FSM_dct_8x8_stage_7_0_t149[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t151 = FSM_dct_8x8_stage_7_0_t150[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t152 = i_data_in[FSM_dct_8x8_stage_7_0_t151 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t153 = FSM_dct_8x8_stage_7_0_t148 + FSM_dct_8x8_stage_7_0_t152;
    FSM_dct_8x8_stage_7_0_t154 = FSM_dct_8x8_stage_7_0_t153[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t155 = FSM_dct_8x8_stage_7_0_t143;
    FSM_dct_8x8_stage_7_0_t155[FSM_dct_8x8_stage_7_0_t145 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t154;
    FSM_dct_8x8_stage_7_0_t156 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_7_0_t157 = FSM_dct_8x8_stage_7_0_t156[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t158 = FSM_dct_8x8_stage_7_0_t157[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t159 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_7_0_t160 = FSM_dct_8x8_stage_7_0_t159[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t161 = FSM_dct_8x8_stage_7_0_t160[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t162 = i_data_in[FSM_dct_8x8_stage_7_0_t161 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t163 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_7_0_t164 = FSM_dct_8x8_stage_7_0_t163[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t165 = FSM_dct_8x8_stage_7_0_t164[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t166 = i_data_in[FSM_dct_8x8_stage_7_0_t165 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t167 = FSM_dct_8x8_stage_7_0_t162 + FSM_dct_8x8_stage_7_0_t166;
    FSM_dct_8x8_stage_7_0_t168 = FSM_dct_8x8_stage_7_0_t167[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t169 = FSM_dct_8x8_stage_7_0_t155;
    FSM_dct_8x8_stage_7_0_t169[FSM_dct_8x8_stage_7_0_t158 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t168;
    FSM_dct_8x8_stage_7_0_t170 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_7_0_t171 = FSM_dct_8x8_stage_7_0_t170[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t172 = FSM_dct_8x8_stage_7_0_t171[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t173 = FSM_dct_8x8_stage_7_0_t169;
    FSM_dct_8x8_stage_7_0_t173[FSM_dct_8x8_stage_7_0_t172 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t162 - FSM_dct_8x8_stage_7_0_t166;
    FSM_dct_8x8_stage_7_0_t174 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_7_0_t175 = FSM_dct_8x8_stage_7_0_t174[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t176 = FSM_dct_8x8_stage_7_0_t175[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t177 = FSM_dct_8x8_stage_7_0_t173;
    FSM_dct_8x8_stage_7_0_t177[FSM_dct_8x8_stage_7_0_t176 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t148 - FSM_dct_8x8_stage_7_0_t152;
    FSM_dct_8x8_stage_7_0_t178 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_7_0_t179 = FSM_dct_8x8_stage_7_0_t178[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t180 = FSM_dct_8x8_stage_7_0_t179[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t181 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_7_0_t182 = FSM_dct_8x8_stage_7_0_t181[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t183 = FSM_dct_8x8_stage_7_0_t182[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t184 = i_data_in[FSM_dct_8x8_stage_7_0_t183 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t185 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_7_0_t186 = FSM_dct_8x8_stage_7_0_t185[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t187 = FSM_dct_8x8_stage_7_0_t186[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t188 = i_data_in[FSM_dct_8x8_stage_7_0_t187 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t189 = FSM_dct_8x8_stage_7_0_t184 + FSM_dct_8x8_stage_7_0_t188;
    FSM_dct_8x8_stage_7_0_t190 = FSM_dct_8x8_stage_7_0_t189[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t191 = FSM_dct_8x8_stage_7_0_t177;
    FSM_dct_8x8_stage_7_0_t191[FSM_dct_8x8_stage_7_0_t180 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t190;
    FSM_dct_8x8_stage_7_0_t192 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_7_0_t193 = FSM_dct_8x8_stage_7_0_t192[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t194 = FSM_dct_8x8_stage_7_0_t193[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t195 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_7_0_t196 = FSM_dct_8x8_stage_7_0_t195[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t197 = FSM_dct_8x8_stage_7_0_t196[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t198 = i_data_in[FSM_dct_8x8_stage_7_0_t197 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t199 = FSM_dct_8x8_stage_7_0_t188 + FSM_dct_8x8_stage_7_0_t198;
    FSM_dct_8x8_stage_7_0_t200 = FSM_dct_8x8_stage_7_0_t199[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t201 = FSM_dct_8x8_stage_7_0_t191;
    FSM_dct_8x8_stage_7_0_t201[FSM_dct_8x8_stage_7_0_t194 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t200;
    FSM_dct_8x8_stage_7_0_t202 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_7_0_t203 = FSM_dct_8x8_stage_7_0_t202[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t204 = FSM_dct_8x8_stage_7_0_t203[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t205 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_7_0_t206 = FSM_dct_8x8_stage_7_0_t205[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t207 = FSM_dct_8x8_stage_7_0_t206[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t208 = i_data_in[FSM_dct_8x8_stage_7_0_t207 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t209 = FSM_dct_8x8_stage_7_0_t198 + FSM_dct_8x8_stage_7_0_t208;
    FSM_dct_8x8_stage_7_0_t210 = FSM_dct_8x8_stage_7_0_t209[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t211 = FSM_dct_8x8_stage_7_0_t201;
    FSM_dct_8x8_stage_7_0_t211[FSM_dct_8x8_stage_7_0_t204 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t210;
    FSM_dct_8x8_stage_7_0_t212 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_7_0_t213 = FSM_dct_8x8_stage_7_0_t212[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t214 = FSM_dct_8x8_stage_7_0_t213[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t215 = FSM_dct_8x8_stage_7_0_t211;
    FSM_dct_8x8_stage_7_0_t215[FSM_dct_8x8_stage_7_0_t214 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t208;
    FSM_dct_8x8_stage_7_0_t216 = 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_7_0_t217 = FSM_dct_8x8_stage_7_0_t216[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t218 = 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_7_0_t219 = FSM_dct_8x8_stage_7_0_t218[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t220 = i_data_in[FSM_dct_8x8_stage_7_0_t219 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t221 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_7_0_t222 = FSM_dct_8x8_stage_7_0_t221[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t223 = FSM_dct_8x8_stage_7_0_t222[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t224 = i_data_in[FSM_dct_8x8_stage_7_0_t223 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t225 = FSM_dct_8x8_stage_7_0_t220 + FSM_dct_8x8_stage_7_0_t224;
    FSM_dct_8x8_stage_7_0_t226 = FSM_dct_8x8_stage_7_0_t225[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t227 = FSM_dct_8x8_stage_7_0_t215;
    FSM_dct_8x8_stage_7_0_t227[FSM_dct_8x8_stage_7_0_t217 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t226;
    FSM_dct_8x8_stage_7_0_t228 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_7_0_t229 = FSM_dct_8x8_stage_7_0_t228[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t230 = FSM_dct_8x8_stage_7_0_t229[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t231 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_7_0_t232 = FSM_dct_8x8_stage_7_0_t231[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t233 = FSM_dct_8x8_stage_7_0_t232[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t234 = i_data_in[FSM_dct_8x8_stage_7_0_t233 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t235 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_7_0_t236 = FSM_dct_8x8_stage_7_0_t235[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t237 = FSM_dct_8x8_stage_7_0_t236[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t238 = i_data_in[FSM_dct_8x8_stage_7_0_t237 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t239 = FSM_dct_8x8_stage_7_0_t234 + FSM_dct_8x8_stage_7_0_t238;
    FSM_dct_8x8_stage_7_0_t240 = FSM_dct_8x8_stage_7_0_t239[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t241 = FSM_dct_8x8_stage_7_0_t227;
    FSM_dct_8x8_stage_7_0_t241[FSM_dct_8x8_stage_7_0_t230 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t240;
    FSM_dct_8x8_stage_7_0_t242 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_7_0_t243 = FSM_dct_8x8_stage_7_0_t242[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t244 = FSM_dct_8x8_stage_7_0_t243[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t245 = FSM_dct_8x8_stage_7_0_t241;
    FSM_dct_8x8_stage_7_0_t245[FSM_dct_8x8_stage_7_0_t244 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t234 - FSM_dct_8x8_stage_7_0_t238;
    FSM_dct_8x8_stage_7_0_t246 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_7_0_t247 = FSM_dct_8x8_stage_7_0_t246[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t248 = FSM_dct_8x8_stage_7_0_t247[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t249 = FSM_dct_8x8_stage_7_0_t245;
    FSM_dct_8x8_stage_7_0_t249[FSM_dct_8x8_stage_7_0_t248 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t220 - FSM_dct_8x8_stage_7_0_t224;
    FSM_dct_8x8_stage_7_0_t250 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_7_0_t251 = FSM_dct_8x8_stage_7_0_t250[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t252 = FSM_dct_8x8_stage_7_0_t251[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t253 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_7_0_t254 = FSM_dct_8x8_stage_7_0_t253[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t255 = FSM_dct_8x8_stage_7_0_t254[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t256 = i_data_in[FSM_dct_8x8_stage_7_0_t255 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t257 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_7_0_t258 = FSM_dct_8x8_stage_7_0_t257[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t259 = FSM_dct_8x8_stage_7_0_t258[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t260 = i_data_in[FSM_dct_8x8_stage_7_0_t259 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t261 = FSM_dct_8x8_stage_7_0_t256 + FSM_dct_8x8_stage_7_0_t260;
    FSM_dct_8x8_stage_7_0_t262 = FSM_dct_8x8_stage_7_0_t261[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t263 = FSM_dct_8x8_stage_7_0_t249;
    FSM_dct_8x8_stage_7_0_t263[FSM_dct_8x8_stage_7_0_t252 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t262;
    FSM_dct_8x8_stage_7_0_t264 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_7_0_t265 = FSM_dct_8x8_stage_7_0_t264[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t266 = FSM_dct_8x8_stage_7_0_t265[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t267 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_7_0_t268 = FSM_dct_8x8_stage_7_0_t267[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t269 = FSM_dct_8x8_stage_7_0_t268[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t270 = i_data_in[FSM_dct_8x8_stage_7_0_t269 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t271 = FSM_dct_8x8_stage_7_0_t260 + FSM_dct_8x8_stage_7_0_t270;
    FSM_dct_8x8_stage_7_0_t272 = FSM_dct_8x8_stage_7_0_t271[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t273 = FSM_dct_8x8_stage_7_0_t263;
    FSM_dct_8x8_stage_7_0_t273[FSM_dct_8x8_stage_7_0_t266 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t272;
    FSM_dct_8x8_stage_7_0_t274 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_7_0_t275 = FSM_dct_8x8_stage_7_0_t274[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t276 = FSM_dct_8x8_stage_7_0_t275[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t277 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_7_0_t278 = FSM_dct_8x8_stage_7_0_t277[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t279 = FSM_dct_8x8_stage_7_0_t278[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t280 = i_data_in[FSM_dct_8x8_stage_7_0_t279 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t281 = FSM_dct_8x8_stage_7_0_t270 + FSM_dct_8x8_stage_7_0_t280;
    FSM_dct_8x8_stage_7_0_t282 = FSM_dct_8x8_stage_7_0_t281[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t283 = FSM_dct_8x8_stage_7_0_t273;
    FSM_dct_8x8_stage_7_0_t283[FSM_dct_8x8_stage_7_0_t276 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t282;
    FSM_dct_8x8_stage_7_0_t284 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_7_0_t285 = FSM_dct_8x8_stage_7_0_t284[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t286 = FSM_dct_8x8_stage_7_0_t285[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t287 = FSM_dct_8x8_stage_7_0_t283;
    FSM_dct_8x8_stage_7_0_t287[FSM_dct_8x8_stage_7_0_t286 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t280;
    FSM_dct_8x8_stage_7_0_t288 = 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_7_0_t289 = FSM_dct_8x8_stage_7_0_t288[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t290 = 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_7_0_t291 = FSM_dct_8x8_stage_7_0_t290[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t292 = i_data_in[FSM_dct_8x8_stage_7_0_t291 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t293 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_7_0_t294 = FSM_dct_8x8_stage_7_0_t293[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t295 = FSM_dct_8x8_stage_7_0_t294[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t296 = i_data_in[FSM_dct_8x8_stage_7_0_t295 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t297 = FSM_dct_8x8_stage_7_0_t292 + FSM_dct_8x8_stage_7_0_t296;
    FSM_dct_8x8_stage_7_0_t298 = FSM_dct_8x8_stage_7_0_t297[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t299 = FSM_dct_8x8_stage_7_0_t287;
    FSM_dct_8x8_stage_7_0_t299[FSM_dct_8x8_stage_7_0_t289 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t298;
    FSM_dct_8x8_stage_7_0_t300 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_7_0_t301 = FSM_dct_8x8_stage_7_0_t300[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t302 = FSM_dct_8x8_stage_7_0_t301[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t303 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_7_0_t304 = FSM_dct_8x8_stage_7_0_t303[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t305 = FSM_dct_8x8_stage_7_0_t304[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t306 = i_data_in[FSM_dct_8x8_stage_7_0_t305 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t307 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_7_0_t308 = FSM_dct_8x8_stage_7_0_t307[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t309 = FSM_dct_8x8_stage_7_0_t308[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t310 = i_data_in[FSM_dct_8x8_stage_7_0_t309 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t311 = FSM_dct_8x8_stage_7_0_t306 + FSM_dct_8x8_stage_7_0_t310;
    FSM_dct_8x8_stage_7_0_t312 = FSM_dct_8x8_stage_7_0_t311[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t313 = FSM_dct_8x8_stage_7_0_t299;
    FSM_dct_8x8_stage_7_0_t313[FSM_dct_8x8_stage_7_0_t302 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t312;
    FSM_dct_8x8_stage_7_0_t314 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_7_0_t315 = FSM_dct_8x8_stage_7_0_t314[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t316 = FSM_dct_8x8_stage_7_0_t315[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t317 = FSM_dct_8x8_stage_7_0_t313;
    FSM_dct_8x8_stage_7_0_t317[FSM_dct_8x8_stage_7_0_t316 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t306 - FSM_dct_8x8_stage_7_0_t310;
    FSM_dct_8x8_stage_7_0_t318 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_7_0_t319 = FSM_dct_8x8_stage_7_0_t318[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t320 = FSM_dct_8x8_stage_7_0_t319[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t321 = FSM_dct_8x8_stage_7_0_t317;
    FSM_dct_8x8_stage_7_0_t321[FSM_dct_8x8_stage_7_0_t320 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t292 - FSM_dct_8x8_stage_7_0_t296;
    FSM_dct_8x8_stage_7_0_t322 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_7_0_t323 = FSM_dct_8x8_stage_7_0_t322[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t324 = FSM_dct_8x8_stage_7_0_t323[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t325 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_7_0_t326 = FSM_dct_8x8_stage_7_0_t325[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t327 = FSM_dct_8x8_stage_7_0_t326[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t328 = i_data_in[FSM_dct_8x8_stage_7_0_t327 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t329 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_7_0_t330 = FSM_dct_8x8_stage_7_0_t329[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t331 = FSM_dct_8x8_stage_7_0_t330[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t332 = i_data_in[FSM_dct_8x8_stage_7_0_t331 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t333 = FSM_dct_8x8_stage_7_0_t328 + FSM_dct_8x8_stage_7_0_t332;
    FSM_dct_8x8_stage_7_0_t334 = FSM_dct_8x8_stage_7_0_t333[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t335 = FSM_dct_8x8_stage_7_0_t321;
    FSM_dct_8x8_stage_7_0_t335[FSM_dct_8x8_stage_7_0_t324 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t334;
    FSM_dct_8x8_stage_7_0_t336 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_7_0_t337 = FSM_dct_8x8_stage_7_0_t336[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t338 = FSM_dct_8x8_stage_7_0_t337[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t339 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_7_0_t340 = FSM_dct_8x8_stage_7_0_t339[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t341 = FSM_dct_8x8_stage_7_0_t340[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t342 = i_data_in[FSM_dct_8x8_stage_7_0_t341 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t343 = FSM_dct_8x8_stage_7_0_t332 + FSM_dct_8x8_stage_7_0_t342;
    FSM_dct_8x8_stage_7_0_t344 = FSM_dct_8x8_stage_7_0_t343[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t345 = FSM_dct_8x8_stage_7_0_t335;
    FSM_dct_8x8_stage_7_0_t345[FSM_dct_8x8_stage_7_0_t338 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t344;
    FSM_dct_8x8_stage_7_0_t346 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_7_0_t347 = FSM_dct_8x8_stage_7_0_t346[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t348 = FSM_dct_8x8_stage_7_0_t347[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t349 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_7_0_t350 = FSM_dct_8x8_stage_7_0_t349[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t351 = FSM_dct_8x8_stage_7_0_t350[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t352 = i_data_in[FSM_dct_8x8_stage_7_0_t351 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t353 = FSM_dct_8x8_stage_7_0_t342 + FSM_dct_8x8_stage_7_0_t352;
    FSM_dct_8x8_stage_7_0_t354 = FSM_dct_8x8_stage_7_0_t353[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t355 = FSM_dct_8x8_stage_7_0_t345;
    FSM_dct_8x8_stage_7_0_t355[FSM_dct_8x8_stage_7_0_t348 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t354;
    FSM_dct_8x8_stage_7_0_t356 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_7_0_t357 = FSM_dct_8x8_stage_7_0_t356[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t358 = FSM_dct_8x8_stage_7_0_t357[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t359 = FSM_dct_8x8_stage_7_0_t355;
    FSM_dct_8x8_stage_7_0_t359[FSM_dct_8x8_stage_7_0_t358 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t352;
    FSM_dct_8x8_stage_7_0_t360 = 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_7_0_t361 = FSM_dct_8x8_stage_7_0_t360[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t362 = 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_7_0_t363 = FSM_dct_8x8_stage_7_0_t362[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t364 = i_data_in[FSM_dct_8x8_stage_7_0_t363 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t365 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_7_0_t366 = FSM_dct_8x8_stage_7_0_t365[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t367 = FSM_dct_8x8_stage_7_0_t366[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t368 = i_data_in[FSM_dct_8x8_stage_7_0_t367 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t369 = FSM_dct_8x8_stage_7_0_t364 + FSM_dct_8x8_stage_7_0_t368;
    FSM_dct_8x8_stage_7_0_t370 = FSM_dct_8x8_stage_7_0_t369[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t371 = FSM_dct_8x8_stage_7_0_t359;
    FSM_dct_8x8_stage_7_0_t371[FSM_dct_8x8_stage_7_0_t361 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t370;
    FSM_dct_8x8_stage_7_0_t372 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_7_0_t373 = FSM_dct_8x8_stage_7_0_t372[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t374 = FSM_dct_8x8_stage_7_0_t373[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t375 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_7_0_t376 = FSM_dct_8x8_stage_7_0_t375[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t377 = FSM_dct_8x8_stage_7_0_t376[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t378 = i_data_in[FSM_dct_8x8_stage_7_0_t377 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t379 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_7_0_t380 = FSM_dct_8x8_stage_7_0_t379[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t381 = FSM_dct_8x8_stage_7_0_t380[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t382 = i_data_in[FSM_dct_8x8_stage_7_0_t381 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t383 = FSM_dct_8x8_stage_7_0_t378 + FSM_dct_8x8_stage_7_0_t382;
    FSM_dct_8x8_stage_7_0_t384 = FSM_dct_8x8_stage_7_0_t383[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t385 = FSM_dct_8x8_stage_7_0_t371;
    FSM_dct_8x8_stage_7_0_t385[FSM_dct_8x8_stage_7_0_t374 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t384;
    FSM_dct_8x8_stage_7_0_t386 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_7_0_t387 = FSM_dct_8x8_stage_7_0_t386[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t388 = FSM_dct_8x8_stage_7_0_t387[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t389 = FSM_dct_8x8_stage_7_0_t385;
    FSM_dct_8x8_stage_7_0_t389[FSM_dct_8x8_stage_7_0_t388 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t378 - FSM_dct_8x8_stage_7_0_t382;
    FSM_dct_8x8_stage_7_0_t390 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_7_0_t391 = FSM_dct_8x8_stage_7_0_t390[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t392 = FSM_dct_8x8_stage_7_0_t391[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t393 = FSM_dct_8x8_stage_7_0_t389;
    FSM_dct_8x8_stage_7_0_t393[FSM_dct_8x8_stage_7_0_t392 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t364 - FSM_dct_8x8_stage_7_0_t368;
    FSM_dct_8x8_stage_7_0_t394 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_7_0_t395 = FSM_dct_8x8_stage_7_0_t394[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t396 = FSM_dct_8x8_stage_7_0_t395[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t397 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_7_0_t398 = FSM_dct_8x8_stage_7_0_t397[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t399 = FSM_dct_8x8_stage_7_0_t398[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t400 = i_data_in[FSM_dct_8x8_stage_7_0_t399 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t401 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_7_0_t402 = FSM_dct_8x8_stage_7_0_t401[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t403 = FSM_dct_8x8_stage_7_0_t402[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t404 = i_data_in[FSM_dct_8x8_stage_7_0_t403 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t405 = FSM_dct_8x8_stage_7_0_t400 + FSM_dct_8x8_stage_7_0_t404;
    FSM_dct_8x8_stage_7_0_t406 = FSM_dct_8x8_stage_7_0_t405[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t407 = FSM_dct_8x8_stage_7_0_t393;
    FSM_dct_8x8_stage_7_0_t407[FSM_dct_8x8_stage_7_0_t396 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t406;
    FSM_dct_8x8_stage_7_0_t408 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_7_0_t409 = FSM_dct_8x8_stage_7_0_t408[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t410 = FSM_dct_8x8_stage_7_0_t409[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t411 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_7_0_t412 = FSM_dct_8x8_stage_7_0_t411[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t413 = FSM_dct_8x8_stage_7_0_t412[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t414 = i_data_in[FSM_dct_8x8_stage_7_0_t413 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t415 = FSM_dct_8x8_stage_7_0_t404 + FSM_dct_8x8_stage_7_0_t414;
    FSM_dct_8x8_stage_7_0_t416 = FSM_dct_8x8_stage_7_0_t415[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t417 = FSM_dct_8x8_stage_7_0_t407;
    FSM_dct_8x8_stage_7_0_t417[FSM_dct_8x8_stage_7_0_t410 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t416;
    FSM_dct_8x8_stage_7_0_t418 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_7_0_t419 = FSM_dct_8x8_stage_7_0_t418[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t420 = FSM_dct_8x8_stage_7_0_t419[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t421 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_7_0_t422 = FSM_dct_8x8_stage_7_0_t421[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t423 = FSM_dct_8x8_stage_7_0_t422[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t424 = i_data_in[FSM_dct_8x8_stage_7_0_t423 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t425 = FSM_dct_8x8_stage_7_0_t414 + FSM_dct_8x8_stage_7_0_t424;
    FSM_dct_8x8_stage_7_0_t426 = FSM_dct_8x8_stage_7_0_t425[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t427 = FSM_dct_8x8_stage_7_0_t417;
    FSM_dct_8x8_stage_7_0_t427[FSM_dct_8x8_stage_7_0_t420 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t426;
    FSM_dct_8x8_stage_7_0_t428 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_7_0_t429 = FSM_dct_8x8_stage_7_0_t428[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t430 = FSM_dct_8x8_stage_7_0_t429[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t431 = FSM_dct_8x8_stage_7_0_t427;
    FSM_dct_8x8_stage_7_0_t431[FSM_dct_8x8_stage_7_0_t430 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t424;
    FSM_dct_8x8_stage_7_0_t432 = 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_7_0_t433 = FSM_dct_8x8_stage_7_0_t432[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t434 = 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_7_0_t435 = FSM_dct_8x8_stage_7_0_t434[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t436 = i_data_in[FSM_dct_8x8_stage_7_0_t435 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t437 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_7_0_t438 = FSM_dct_8x8_stage_7_0_t437[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t439 = FSM_dct_8x8_stage_7_0_t438[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t440 = i_data_in[FSM_dct_8x8_stage_7_0_t439 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t441 = FSM_dct_8x8_stage_7_0_t436 + FSM_dct_8x8_stage_7_0_t440;
    FSM_dct_8x8_stage_7_0_t442 = FSM_dct_8x8_stage_7_0_t441[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t443 = FSM_dct_8x8_stage_7_0_t431;
    FSM_dct_8x8_stage_7_0_t443[FSM_dct_8x8_stage_7_0_t433 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t442;
    FSM_dct_8x8_stage_7_0_t444 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_7_0_t445 = FSM_dct_8x8_stage_7_0_t444[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t446 = FSM_dct_8x8_stage_7_0_t445[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t447 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_7_0_t448 = FSM_dct_8x8_stage_7_0_t447[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t449 = FSM_dct_8x8_stage_7_0_t448[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t450 = i_data_in[FSM_dct_8x8_stage_7_0_t449 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t451 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_7_0_t452 = FSM_dct_8x8_stage_7_0_t451[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t453 = FSM_dct_8x8_stage_7_0_t452[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t454 = i_data_in[FSM_dct_8x8_stage_7_0_t453 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t455 = FSM_dct_8x8_stage_7_0_t450 + FSM_dct_8x8_stage_7_0_t454;
    FSM_dct_8x8_stage_7_0_t456 = FSM_dct_8x8_stage_7_0_t455[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t457 = FSM_dct_8x8_stage_7_0_t443;
    FSM_dct_8x8_stage_7_0_t457[FSM_dct_8x8_stage_7_0_t446 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t456;
    FSM_dct_8x8_stage_7_0_t458 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_7_0_t459 = FSM_dct_8x8_stage_7_0_t458[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t460 = FSM_dct_8x8_stage_7_0_t459[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t461 = FSM_dct_8x8_stage_7_0_t457;
    FSM_dct_8x8_stage_7_0_t461[FSM_dct_8x8_stage_7_0_t460 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t450 - FSM_dct_8x8_stage_7_0_t454;
    FSM_dct_8x8_stage_7_0_t462 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_7_0_t463 = FSM_dct_8x8_stage_7_0_t462[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t464 = FSM_dct_8x8_stage_7_0_t463[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t465 = FSM_dct_8x8_stage_7_0_t461;
    FSM_dct_8x8_stage_7_0_t465[FSM_dct_8x8_stage_7_0_t464 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t436 - FSM_dct_8x8_stage_7_0_t440;
    FSM_dct_8x8_stage_7_0_t466 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_7_0_t467 = FSM_dct_8x8_stage_7_0_t466[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t468 = FSM_dct_8x8_stage_7_0_t467[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t469 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_7_0_t470 = FSM_dct_8x8_stage_7_0_t469[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t471 = FSM_dct_8x8_stage_7_0_t470[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t472 = i_data_in[FSM_dct_8x8_stage_7_0_t471 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t473 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_7_0_t474 = FSM_dct_8x8_stage_7_0_t473[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t475 = FSM_dct_8x8_stage_7_0_t474[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t476 = i_data_in[FSM_dct_8x8_stage_7_0_t475 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t477 = FSM_dct_8x8_stage_7_0_t472 + FSM_dct_8x8_stage_7_0_t476;
    FSM_dct_8x8_stage_7_0_t478 = FSM_dct_8x8_stage_7_0_t477[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t479 = FSM_dct_8x8_stage_7_0_t465;
    FSM_dct_8x8_stage_7_0_t479[FSM_dct_8x8_stage_7_0_t468 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t478;
    FSM_dct_8x8_stage_7_0_t480 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_7_0_t481 = FSM_dct_8x8_stage_7_0_t480[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t482 = FSM_dct_8x8_stage_7_0_t481[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t483 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_7_0_t484 = FSM_dct_8x8_stage_7_0_t483[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t485 = FSM_dct_8x8_stage_7_0_t484[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t486 = i_data_in[FSM_dct_8x8_stage_7_0_t485 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t487 = FSM_dct_8x8_stage_7_0_t476 + FSM_dct_8x8_stage_7_0_t486;
    FSM_dct_8x8_stage_7_0_t488 = FSM_dct_8x8_stage_7_0_t487[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t489 = FSM_dct_8x8_stage_7_0_t479;
    FSM_dct_8x8_stage_7_0_t489[FSM_dct_8x8_stage_7_0_t482 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t488;
    FSM_dct_8x8_stage_7_0_t490 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_7_0_t491 = FSM_dct_8x8_stage_7_0_t490[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t492 = FSM_dct_8x8_stage_7_0_t491[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t493 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_7_0_t494 = FSM_dct_8x8_stage_7_0_t493[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t495 = FSM_dct_8x8_stage_7_0_t494[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t496 = i_data_in[FSM_dct_8x8_stage_7_0_t495 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t497 = FSM_dct_8x8_stage_7_0_t486 + FSM_dct_8x8_stage_7_0_t496;
    FSM_dct_8x8_stage_7_0_t498 = FSM_dct_8x8_stage_7_0_t497[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t499 = FSM_dct_8x8_stage_7_0_t489;
    FSM_dct_8x8_stage_7_0_t499[FSM_dct_8x8_stage_7_0_t492 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t498;
    FSM_dct_8x8_stage_7_0_t500 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_7_0_t501 = FSM_dct_8x8_stage_7_0_t500[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t502 = FSM_dct_8x8_stage_7_0_t501[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t503 = FSM_dct_8x8_stage_7_0_t499;
    FSM_dct_8x8_stage_7_0_t503[FSM_dct_8x8_stage_7_0_t502 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t496;
    FSM_dct_8x8_stage_7_0_t504 = 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_7_0_t505 = FSM_dct_8x8_stage_7_0_t504[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t506 = 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_7_0_t507 = FSM_dct_8x8_stage_7_0_t506[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t508 = i_data_in[FSM_dct_8x8_stage_7_0_t507 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t509 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_7_0_t510 = FSM_dct_8x8_stage_7_0_t509[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t511 = FSM_dct_8x8_stage_7_0_t510[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t512 = i_data_in[FSM_dct_8x8_stage_7_0_t511 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t513 = FSM_dct_8x8_stage_7_0_t508 + FSM_dct_8x8_stage_7_0_t512;
    FSM_dct_8x8_stage_7_0_t514 = FSM_dct_8x8_stage_7_0_t513[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t515 = FSM_dct_8x8_stage_7_0_t503;
    FSM_dct_8x8_stage_7_0_t515[FSM_dct_8x8_stage_7_0_t505 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t514;
    FSM_dct_8x8_stage_7_0_t516 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_7_0_t517 = FSM_dct_8x8_stage_7_0_t516[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t518 = FSM_dct_8x8_stage_7_0_t517[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t519 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_7_0_t520 = FSM_dct_8x8_stage_7_0_t519[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t521 = FSM_dct_8x8_stage_7_0_t520[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t522 = i_data_in[FSM_dct_8x8_stage_7_0_t521 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t523 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_7_0_t524 = FSM_dct_8x8_stage_7_0_t523[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t525 = FSM_dct_8x8_stage_7_0_t524[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t526 = i_data_in[FSM_dct_8x8_stage_7_0_t525 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t527 = FSM_dct_8x8_stage_7_0_t522 + FSM_dct_8x8_stage_7_0_t526;
    FSM_dct_8x8_stage_7_0_t528 = FSM_dct_8x8_stage_7_0_t527[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t529 = FSM_dct_8x8_stage_7_0_t515;
    FSM_dct_8x8_stage_7_0_t529[FSM_dct_8x8_stage_7_0_t518 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t528;
    FSM_dct_8x8_stage_7_0_t530 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_7_0_t531 = FSM_dct_8x8_stage_7_0_t530[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t532 = FSM_dct_8x8_stage_7_0_t531[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t533 = FSM_dct_8x8_stage_7_0_t529;
    FSM_dct_8x8_stage_7_0_t533[FSM_dct_8x8_stage_7_0_t532 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t522 - FSM_dct_8x8_stage_7_0_t526;
    FSM_dct_8x8_stage_7_0_t534 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_7_0_t535 = FSM_dct_8x8_stage_7_0_t534[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t536 = FSM_dct_8x8_stage_7_0_t535[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t537 = FSM_dct_8x8_stage_7_0_t533;
    FSM_dct_8x8_stage_7_0_t537[FSM_dct_8x8_stage_7_0_t536 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t508 - FSM_dct_8x8_stage_7_0_t512;
    FSM_dct_8x8_stage_7_0_t538 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_7_0_t539 = FSM_dct_8x8_stage_7_0_t538[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t540 = FSM_dct_8x8_stage_7_0_t539[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t541 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_7_0_t542 = FSM_dct_8x8_stage_7_0_t541[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t543 = FSM_dct_8x8_stage_7_0_t542[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t544 = i_data_in[FSM_dct_8x8_stage_7_0_t543 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t545 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_7_0_t546 = FSM_dct_8x8_stage_7_0_t545[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t547 = FSM_dct_8x8_stage_7_0_t546[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t548 = i_data_in[FSM_dct_8x8_stage_7_0_t547 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t549 = FSM_dct_8x8_stage_7_0_t544 + FSM_dct_8x8_stage_7_0_t548;
    FSM_dct_8x8_stage_7_0_t550 = FSM_dct_8x8_stage_7_0_t549[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t551 = FSM_dct_8x8_stage_7_0_t537;
    FSM_dct_8x8_stage_7_0_t551[FSM_dct_8x8_stage_7_0_t540 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t550;
    FSM_dct_8x8_stage_7_0_t552 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_7_0_t553 = FSM_dct_8x8_stage_7_0_t552[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t554 = FSM_dct_8x8_stage_7_0_t553[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t555 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_7_0_t556 = FSM_dct_8x8_stage_7_0_t555[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t557 = FSM_dct_8x8_stage_7_0_t556[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t558 = i_data_in[FSM_dct_8x8_stage_7_0_t557 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t559 = FSM_dct_8x8_stage_7_0_t548 + FSM_dct_8x8_stage_7_0_t558;
    FSM_dct_8x8_stage_7_0_t560 = FSM_dct_8x8_stage_7_0_t559[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t561 = FSM_dct_8x8_stage_7_0_t551;
    FSM_dct_8x8_stage_7_0_t561[FSM_dct_8x8_stage_7_0_t554 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t560;
    FSM_dct_8x8_stage_7_0_t562 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_7_0_t563 = FSM_dct_8x8_stage_7_0_t562[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t564 = FSM_dct_8x8_stage_7_0_t563[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t565 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_7_0_t566 = FSM_dct_8x8_stage_7_0_t565[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t567 = FSM_dct_8x8_stage_7_0_t566[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t568 = i_data_in[FSM_dct_8x8_stage_7_0_t567 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t569 = FSM_dct_8x8_stage_7_0_t558 + FSM_dct_8x8_stage_7_0_t568;
    FSM_dct_8x8_stage_7_0_t570 = FSM_dct_8x8_stage_7_0_t569[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t571 = FSM_dct_8x8_stage_7_0_t561;
    FSM_dct_8x8_stage_7_0_t571[FSM_dct_8x8_stage_7_0_t564 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t570;
    FSM_dct_8x8_stage_7_0_t572 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_7_0_t573 = FSM_dct_8x8_stage_7_0_t572[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t574 = FSM_dct_8x8_stage_7_0_t573[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t575 = FSM_dct_8x8_stage_7_0_t571;
    FSM_dct_8x8_stage_7_0_t575[FSM_dct_8x8_stage_7_0_t574 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t568;
end

always @* begin
    FSM_dct_8x8_stage_7_0_t0 = 32'b0;
    FSM_dct_8x8_stage_7_0_t1 = FSM_dct_8x8_stage_7_0_t0[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t2 = 32'b0;
    FSM_dct_8x8_stage_7_0_t3 = FSM_dct_8x8_stage_7_0_t2[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t4 = i_data_in[FSM_dct_8x8_stage_7_0_t3 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t5 = 32'b00000000000000000000000000011000 + 32'b0;
    FSM_dct_8x8_stage_7_0_t6 = FSM_dct_8x8_stage_7_0_t5[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t7 = FSM_dct_8x8_stage_7_0_t6[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t8 = i_data_in[FSM_dct_8x8_stage_7_0_t7 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t9 = FSM_dct_8x8_stage_7_0_t4 + FSM_dct_8x8_stage_7_0_t8;
    FSM_dct_8x8_stage_7_0_t10 = FSM_dct_8x8_stage_7_0_t9[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t11 = 2048'b0;
    FSM_dct_8x8_stage_7_0_t11[FSM_dct_8x8_stage_7_0_t1 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t10;
    FSM_dct_8x8_stage_7_0_t12 = 32'b00000000000000000000000000001000 + 32'b0;
    FSM_dct_8x8_stage_7_0_t13 = FSM_dct_8x8_stage_7_0_t12[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t14 = FSM_dct_8x8_stage_7_0_t13[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t15 = 32'b00000000000000000000000000001000 + 32'b0;
    FSM_dct_8x8_stage_7_0_t16 = FSM_dct_8x8_stage_7_0_t15[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t17 = FSM_dct_8x8_stage_7_0_t16[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t18 = i_data_in[FSM_dct_8x8_stage_7_0_t17 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t19 = 32'b00000000000000000000000000010000 + 32'b0;
    FSM_dct_8x8_stage_7_0_t20 = FSM_dct_8x8_stage_7_0_t19[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t21 = FSM_dct_8x8_stage_7_0_t20[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t22 = i_data_in[FSM_dct_8x8_stage_7_0_t21 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t23 = FSM_dct_8x8_stage_7_0_t18 + FSM_dct_8x8_stage_7_0_t22;
    FSM_dct_8x8_stage_7_0_t24 = FSM_dct_8x8_stage_7_0_t23[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t25 = FSM_dct_8x8_stage_7_0_t11;
    FSM_dct_8x8_stage_7_0_t25[FSM_dct_8x8_stage_7_0_t14 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t24;
    FSM_dct_8x8_stage_7_0_t26 = 32'b00000000000000000000000000010000 + 32'b0;
    FSM_dct_8x8_stage_7_0_t27 = FSM_dct_8x8_stage_7_0_t26[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t28 = FSM_dct_8x8_stage_7_0_t27[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t29 = FSM_dct_8x8_stage_7_0_t25;
    FSM_dct_8x8_stage_7_0_t29[FSM_dct_8x8_stage_7_0_t28 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t18 - FSM_dct_8x8_stage_7_0_t22;
    FSM_dct_8x8_stage_7_0_t30 = 32'b00000000000000000000000000011000 + 32'b0;
    FSM_dct_8x8_stage_7_0_t31 = FSM_dct_8x8_stage_7_0_t30[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t32 = FSM_dct_8x8_stage_7_0_t31[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t33 = FSM_dct_8x8_stage_7_0_t29;
    FSM_dct_8x8_stage_7_0_t33[FSM_dct_8x8_stage_7_0_t32 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t4 - FSM_dct_8x8_stage_7_0_t8;
    FSM_dct_8x8_stage_7_0_t34 = 32'b00000000000000000000000000100000 + 32'b0;
    FSM_dct_8x8_stage_7_0_t35 = FSM_dct_8x8_stage_7_0_t34[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t36 = FSM_dct_8x8_stage_7_0_t35[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t37 = 32'b00000000000000000000000000100000 + 32'b0;
    FSM_dct_8x8_stage_7_0_t38 = FSM_dct_8x8_stage_7_0_t37[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t39 = FSM_dct_8x8_stage_7_0_t38[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t40 = i_data_in[FSM_dct_8x8_stage_7_0_t39 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t41 = 32'b00000000000000000000000000101000 + 32'b0;
    FSM_dct_8x8_stage_7_0_t42 = FSM_dct_8x8_stage_7_0_t41[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t43 = FSM_dct_8x8_stage_7_0_t42[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t44 = i_data_in[FSM_dct_8x8_stage_7_0_t43 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t45 = FSM_dct_8x8_stage_7_0_t40 + FSM_dct_8x8_stage_7_0_t44;
    FSM_dct_8x8_stage_7_0_t46 = FSM_dct_8x8_stage_7_0_t45[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t47 = FSM_dct_8x8_stage_7_0_t33;
    FSM_dct_8x8_stage_7_0_t47[FSM_dct_8x8_stage_7_0_t36 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t46;
    FSM_dct_8x8_stage_7_0_t48 = 32'b00000000000000000000000000101000 + 32'b0;
    FSM_dct_8x8_stage_7_0_t49 = FSM_dct_8x8_stage_7_0_t48[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t50 = FSM_dct_8x8_stage_7_0_t49[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t51 = 32'b00000000000000000000000000110000 + 32'b0;
    FSM_dct_8x8_stage_7_0_t52 = FSM_dct_8x8_stage_7_0_t51[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t53 = FSM_dct_8x8_stage_7_0_t52[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t54 = i_data_in[FSM_dct_8x8_stage_7_0_t53 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t55 = FSM_dct_8x8_stage_7_0_t44 + FSM_dct_8x8_stage_7_0_t54;
    FSM_dct_8x8_stage_7_0_t56 = FSM_dct_8x8_stage_7_0_t55[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t57 = FSM_dct_8x8_stage_7_0_t47;
    FSM_dct_8x8_stage_7_0_t57[FSM_dct_8x8_stage_7_0_t50 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t56;
    FSM_dct_8x8_stage_7_0_t58 = 32'b00000000000000000000000000110000 + 32'b0;
    FSM_dct_8x8_stage_7_0_t59 = FSM_dct_8x8_stage_7_0_t58[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t60 = FSM_dct_8x8_stage_7_0_t59[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t61 = 32'b00000000000000000000000000111000 + 32'b0;
    FSM_dct_8x8_stage_7_0_t62 = FSM_dct_8x8_stage_7_0_t61[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t63 = FSM_dct_8x8_stage_7_0_t62[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t64 = i_data_in[FSM_dct_8x8_stage_7_0_t63 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t65 = FSM_dct_8x8_stage_7_0_t54 + FSM_dct_8x8_stage_7_0_t64;
    FSM_dct_8x8_stage_7_0_t66 = FSM_dct_8x8_stage_7_0_t65[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t67 = FSM_dct_8x8_stage_7_0_t57;
    FSM_dct_8x8_stage_7_0_t67[FSM_dct_8x8_stage_7_0_t60 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t66;
    FSM_dct_8x8_stage_7_0_t68 = 32'b00000000000000000000000000111000 + 32'b0;
    FSM_dct_8x8_stage_7_0_t69 = FSM_dct_8x8_stage_7_0_t68[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t70 = FSM_dct_8x8_stage_7_0_t69[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t71 = FSM_dct_8x8_stage_7_0_t67;
    FSM_dct_8x8_stage_7_0_t71[FSM_dct_8x8_stage_7_0_t70 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t64;
    FSM_dct_8x8_stage_7_0_t72 = 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_7_0_t73 = FSM_dct_8x8_stage_7_0_t72[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t74 = 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_7_0_t75 = FSM_dct_8x8_stage_7_0_t74[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t76 = i_data_in[FSM_dct_8x8_stage_7_0_t75 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t77 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_7_0_t78 = FSM_dct_8x8_stage_7_0_t77[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t79 = FSM_dct_8x8_stage_7_0_t78[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t80 = i_data_in[FSM_dct_8x8_stage_7_0_t79 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t81 = FSM_dct_8x8_stage_7_0_t76 + FSM_dct_8x8_stage_7_0_t80;
    FSM_dct_8x8_stage_7_0_t82 = FSM_dct_8x8_stage_7_0_t81[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t83 = FSM_dct_8x8_stage_7_0_t71;
    FSM_dct_8x8_stage_7_0_t83[FSM_dct_8x8_stage_7_0_t73 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t82;
    FSM_dct_8x8_stage_7_0_t84 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_7_0_t85 = FSM_dct_8x8_stage_7_0_t84[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t86 = FSM_dct_8x8_stage_7_0_t85[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t87 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_7_0_t88 = FSM_dct_8x8_stage_7_0_t87[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t89 = FSM_dct_8x8_stage_7_0_t88[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t90 = i_data_in[FSM_dct_8x8_stage_7_0_t89 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t91 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_7_0_t92 = FSM_dct_8x8_stage_7_0_t91[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t93 = FSM_dct_8x8_stage_7_0_t92[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t94 = i_data_in[FSM_dct_8x8_stage_7_0_t93 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t95 = FSM_dct_8x8_stage_7_0_t90 + FSM_dct_8x8_stage_7_0_t94;
    FSM_dct_8x8_stage_7_0_t96 = FSM_dct_8x8_stage_7_0_t95[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t97 = FSM_dct_8x8_stage_7_0_t83;
    FSM_dct_8x8_stage_7_0_t97[FSM_dct_8x8_stage_7_0_t86 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t96;
    FSM_dct_8x8_stage_7_0_t98 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_7_0_t99 = FSM_dct_8x8_stage_7_0_t98[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t100 = FSM_dct_8x8_stage_7_0_t99[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t101 = FSM_dct_8x8_stage_7_0_t97;
    FSM_dct_8x8_stage_7_0_t101[FSM_dct_8x8_stage_7_0_t100 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t90 - FSM_dct_8x8_stage_7_0_t94;
    FSM_dct_8x8_stage_7_0_t102 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_7_0_t103 = FSM_dct_8x8_stage_7_0_t102[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t104 = FSM_dct_8x8_stage_7_0_t103[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t105 = FSM_dct_8x8_stage_7_0_t101;
    FSM_dct_8x8_stage_7_0_t105[FSM_dct_8x8_stage_7_0_t104 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t76 - FSM_dct_8x8_stage_7_0_t80;
    FSM_dct_8x8_stage_7_0_t106 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_7_0_t107 = FSM_dct_8x8_stage_7_0_t106[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t108 = FSM_dct_8x8_stage_7_0_t107[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t109 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_7_0_t110 = FSM_dct_8x8_stage_7_0_t109[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t111 = FSM_dct_8x8_stage_7_0_t110[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t112 = i_data_in[FSM_dct_8x8_stage_7_0_t111 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t113 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_7_0_t114 = FSM_dct_8x8_stage_7_0_t113[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t115 = FSM_dct_8x8_stage_7_0_t114[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t116 = i_data_in[FSM_dct_8x8_stage_7_0_t115 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t117 = FSM_dct_8x8_stage_7_0_t112 + FSM_dct_8x8_stage_7_0_t116;
    FSM_dct_8x8_stage_7_0_t118 = FSM_dct_8x8_stage_7_0_t117[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t119 = FSM_dct_8x8_stage_7_0_t105;
    FSM_dct_8x8_stage_7_0_t119[FSM_dct_8x8_stage_7_0_t108 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t118;
    FSM_dct_8x8_stage_7_0_t120 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_7_0_t121 = FSM_dct_8x8_stage_7_0_t120[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t122 = FSM_dct_8x8_stage_7_0_t121[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t123 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_7_0_t124 = FSM_dct_8x8_stage_7_0_t123[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t125 = FSM_dct_8x8_stage_7_0_t124[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t126 = i_data_in[FSM_dct_8x8_stage_7_0_t125 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t127 = FSM_dct_8x8_stage_7_0_t116 + FSM_dct_8x8_stage_7_0_t126;
    FSM_dct_8x8_stage_7_0_t128 = FSM_dct_8x8_stage_7_0_t127[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t129 = FSM_dct_8x8_stage_7_0_t119;
    FSM_dct_8x8_stage_7_0_t129[FSM_dct_8x8_stage_7_0_t122 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t128;
    FSM_dct_8x8_stage_7_0_t130 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_7_0_t131 = FSM_dct_8x8_stage_7_0_t130[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t132 = FSM_dct_8x8_stage_7_0_t131[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t133 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_7_0_t134 = FSM_dct_8x8_stage_7_0_t133[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t135 = FSM_dct_8x8_stage_7_0_t134[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t136 = i_data_in[FSM_dct_8x8_stage_7_0_t135 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t137 = FSM_dct_8x8_stage_7_0_t126 + FSM_dct_8x8_stage_7_0_t136;
    FSM_dct_8x8_stage_7_0_t138 = FSM_dct_8x8_stage_7_0_t137[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t139 = FSM_dct_8x8_stage_7_0_t129;
    FSM_dct_8x8_stage_7_0_t139[FSM_dct_8x8_stage_7_0_t132 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t138;
    FSM_dct_8x8_stage_7_0_t140 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_7_0_t141 = FSM_dct_8x8_stage_7_0_t140[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t142 = FSM_dct_8x8_stage_7_0_t141[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t143 = FSM_dct_8x8_stage_7_0_t139;
    FSM_dct_8x8_stage_7_0_t143[FSM_dct_8x8_stage_7_0_t142 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t136;
    FSM_dct_8x8_stage_7_0_t144 = 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_7_0_t145 = FSM_dct_8x8_stage_7_0_t144[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t146 = 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_7_0_t147 = FSM_dct_8x8_stage_7_0_t146[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t148 = i_data_in[FSM_dct_8x8_stage_7_0_t147 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t149 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_7_0_t150 = FSM_dct_8x8_stage_7_0_t149[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t151 = FSM_dct_8x8_stage_7_0_t150[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t152 = i_data_in[FSM_dct_8x8_stage_7_0_t151 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t153 = FSM_dct_8x8_stage_7_0_t148 + FSM_dct_8x8_stage_7_0_t152;
    FSM_dct_8x8_stage_7_0_t154 = FSM_dct_8x8_stage_7_0_t153[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t155 = FSM_dct_8x8_stage_7_0_t143;
    FSM_dct_8x8_stage_7_0_t155[FSM_dct_8x8_stage_7_0_t145 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t154;
    FSM_dct_8x8_stage_7_0_t156 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_7_0_t157 = FSM_dct_8x8_stage_7_0_t156[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t158 = FSM_dct_8x8_stage_7_0_t157[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t159 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_7_0_t160 = FSM_dct_8x8_stage_7_0_t159[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t161 = FSM_dct_8x8_stage_7_0_t160[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t162 = i_data_in[FSM_dct_8x8_stage_7_0_t161 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t163 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_7_0_t164 = FSM_dct_8x8_stage_7_0_t163[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t165 = FSM_dct_8x8_stage_7_0_t164[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t166 = i_data_in[FSM_dct_8x8_stage_7_0_t165 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t167 = FSM_dct_8x8_stage_7_0_t162 + FSM_dct_8x8_stage_7_0_t166;
    FSM_dct_8x8_stage_7_0_t168 = FSM_dct_8x8_stage_7_0_t167[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t169 = FSM_dct_8x8_stage_7_0_t155;
    FSM_dct_8x8_stage_7_0_t169[FSM_dct_8x8_stage_7_0_t158 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t168;
    FSM_dct_8x8_stage_7_0_t170 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_7_0_t171 = FSM_dct_8x8_stage_7_0_t170[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t172 = FSM_dct_8x8_stage_7_0_t171[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t173 = FSM_dct_8x8_stage_7_0_t169;
    FSM_dct_8x8_stage_7_0_t173[FSM_dct_8x8_stage_7_0_t172 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t162 - FSM_dct_8x8_stage_7_0_t166;
    FSM_dct_8x8_stage_7_0_t174 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_7_0_t175 = FSM_dct_8x8_stage_7_0_t174[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t176 = FSM_dct_8x8_stage_7_0_t175[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t177 = FSM_dct_8x8_stage_7_0_t173;
    FSM_dct_8x8_stage_7_0_t177[FSM_dct_8x8_stage_7_0_t176 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t148 - FSM_dct_8x8_stage_7_0_t152;
    FSM_dct_8x8_stage_7_0_t178 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_7_0_t179 = FSM_dct_8x8_stage_7_0_t178[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t180 = FSM_dct_8x8_stage_7_0_t179[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t181 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_7_0_t182 = FSM_dct_8x8_stage_7_0_t181[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t183 = FSM_dct_8x8_stage_7_0_t182[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t184 = i_data_in[FSM_dct_8x8_stage_7_0_t183 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t185 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_7_0_t186 = FSM_dct_8x8_stage_7_0_t185[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t187 = FSM_dct_8x8_stage_7_0_t186[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t188 = i_data_in[FSM_dct_8x8_stage_7_0_t187 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t189 = FSM_dct_8x8_stage_7_0_t184 + FSM_dct_8x8_stage_7_0_t188;
    FSM_dct_8x8_stage_7_0_t190 = FSM_dct_8x8_stage_7_0_t189[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t191 = FSM_dct_8x8_stage_7_0_t177;
    FSM_dct_8x8_stage_7_0_t191[FSM_dct_8x8_stage_7_0_t180 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t190;
    FSM_dct_8x8_stage_7_0_t192 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_7_0_t193 = FSM_dct_8x8_stage_7_0_t192[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t194 = FSM_dct_8x8_stage_7_0_t193[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t195 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_7_0_t196 = FSM_dct_8x8_stage_7_0_t195[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t197 = FSM_dct_8x8_stage_7_0_t196[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t198 = i_data_in[FSM_dct_8x8_stage_7_0_t197 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t199 = FSM_dct_8x8_stage_7_0_t188 + FSM_dct_8x8_stage_7_0_t198;
    FSM_dct_8x8_stage_7_0_t200 = FSM_dct_8x8_stage_7_0_t199[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t201 = FSM_dct_8x8_stage_7_0_t191;
    FSM_dct_8x8_stage_7_0_t201[FSM_dct_8x8_stage_7_0_t194 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t200;
    FSM_dct_8x8_stage_7_0_t202 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_7_0_t203 = FSM_dct_8x8_stage_7_0_t202[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t204 = FSM_dct_8x8_stage_7_0_t203[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t205 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_7_0_t206 = FSM_dct_8x8_stage_7_0_t205[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t207 = FSM_dct_8x8_stage_7_0_t206[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t208 = i_data_in[FSM_dct_8x8_stage_7_0_t207 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t209 = FSM_dct_8x8_stage_7_0_t198 + FSM_dct_8x8_stage_7_0_t208;
    FSM_dct_8x8_stage_7_0_t210 = FSM_dct_8x8_stage_7_0_t209[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t211 = FSM_dct_8x8_stage_7_0_t201;
    FSM_dct_8x8_stage_7_0_t211[FSM_dct_8x8_stage_7_0_t204 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t210;
    FSM_dct_8x8_stage_7_0_t212 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_7_0_t213 = FSM_dct_8x8_stage_7_0_t212[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t214 = FSM_dct_8x8_stage_7_0_t213[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t215 = FSM_dct_8x8_stage_7_0_t211;
    FSM_dct_8x8_stage_7_0_t215[FSM_dct_8x8_stage_7_0_t214 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t208;
    FSM_dct_8x8_stage_7_0_t216 = 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_7_0_t217 = FSM_dct_8x8_stage_7_0_t216[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t218 = 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_7_0_t219 = FSM_dct_8x8_stage_7_0_t218[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t220 = i_data_in[FSM_dct_8x8_stage_7_0_t219 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t221 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_7_0_t222 = FSM_dct_8x8_stage_7_0_t221[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t223 = FSM_dct_8x8_stage_7_0_t222[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t224 = i_data_in[FSM_dct_8x8_stage_7_0_t223 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t225 = FSM_dct_8x8_stage_7_0_t220 + FSM_dct_8x8_stage_7_0_t224;
    FSM_dct_8x8_stage_7_0_t226 = FSM_dct_8x8_stage_7_0_t225[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t227 = FSM_dct_8x8_stage_7_0_t215;
    FSM_dct_8x8_stage_7_0_t227[FSM_dct_8x8_stage_7_0_t217 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t226;
    FSM_dct_8x8_stage_7_0_t228 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_7_0_t229 = FSM_dct_8x8_stage_7_0_t228[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t230 = FSM_dct_8x8_stage_7_0_t229[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t231 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_7_0_t232 = FSM_dct_8x8_stage_7_0_t231[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t233 = FSM_dct_8x8_stage_7_0_t232[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t234 = i_data_in[FSM_dct_8x8_stage_7_0_t233 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t235 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_7_0_t236 = FSM_dct_8x8_stage_7_0_t235[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t237 = FSM_dct_8x8_stage_7_0_t236[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t238 = i_data_in[FSM_dct_8x8_stage_7_0_t237 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t239 = FSM_dct_8x8_stage_7_0_t234 + FSM_dct_8x8_stage_7_0_t238;
    FSM_dct_8x8_stage_7_0_t240 = FSM_dct_8x8_stage_7_0_t239[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t241 = FSM_dct_8x8_stage_7_0_t227;
    FSM_dct_8x8_stage_7_0_t241[FSM_dct_8x8_stage_7_0_t230 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t240;
    FSM_dct_8x8_stage_7_0_t242 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_7_0_t243 = FSM_dct_8x8_stage_7_0_t242[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t244 = FSM_dct_8x8_stage_7_0_t243[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t245 = FSM_dct_8x8_stage_7_0_t241;
    FSM_dct_8x8_stage_7_0_t245[FSM_dct_8x8_stage_7_0_t244 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t234 - FSM_dct_8x8_stage_7_0_t238;
    FSM_dct_8x8_stage_7_0_t246 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_7_0_t247 = FSM_dct_8x8_stage_7_0_t246[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t248 = FSM_dct_8x8_stage_7_0_t247[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t249 = FSM_dct_8x8_stage_7_0_t245;
    FSM_dct_8x8_stage_7_0_t249[FSM_dct_8x8_stage_7_0_t248 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t220 - FSM_dct_8x8_stage_7_0_t224;
    FSM_dct_8x8_stage_7_0_t250 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_7_0_t251 = FSM_dct_8x8_stage_7_0_t250[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t252 = FSM_dct_8x8_stage_7_0_t251[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t253 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_7_0_t254 = FSM_dct_8x8_stage_7_0_t253[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t255 = FSM_dct_8x8_stage_7_0_t254[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t256 = i_data_in[FSM_dct_8x8_stage_7_0_t255 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t257 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_7_0_t258 = FSM_dct_8x8_stage_7_0_t257[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t259 = FSM_dct_8x8_stage_7_0_t258[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t260 = i_data_in[FSM_dct_8x8_stage_7_0_t259 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t261 = FSM_dct_8x8_stage_7_0_t256 + FSM_dct_8x8_stage_7_0_t260;
    FSM_dct_8x8_stage_7_0_t262 = FSM_dct_8x8_stage_7_0_t261[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t263 = FSM_dct_8x8_stage_7_0_t249;
    FSM_dct_8x8_stage_7_0_t263[FSM_dct_8x8_stage_7_0_t252 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t262;
    FSM_dct_8x8_stage_7_0_t264 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_7_0_t265 = FSM_dct_8x8_stage_7_0_t264[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t266 = FSM_dct_8x8_stage_7_0_t265[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t267 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_7_0_t268 = FSM_dct_8x8_stage_7_0_t267[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t269 = FSM_dct_8x8_stage_7_0_t268[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t270 = i_data_in[FSM_dct_8x8_stage_7_0_t269 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t271 = FSM_dct_8x8_stage_7_0_t260 + FSM_dct_8x8_stage_7_0_t270;
    FSM_dct_8x8_stage_7_0_t272 = FSM_dct_8x8_stage_7_0_t271[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t273 = FSM_dct_8x8_stage_7_0_t263;
    FSM_dct_8x8_stage_7_0_t273[FSM_dct_8x8_stage_7_0_t266 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t272;
    FSM_dct_8x8_stage_7_0_t274 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_7_0_t275 = FSM_dct_8x8_stage_7_0_t274[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t276 = FSM_dct_8x8_stage_7_0_t275[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t277 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_7_0_t278 = FSM_dct_8x8_stage_7_0_t277[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t279 = FSM_dct_8x8_stage_7_0_t278[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t280 = i_data_in[FSM_dct_8x8_stage_7_0_t279 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t281 = FSM_dct_8x8_stage_7_0_t270 + FSM_dct_8x8_stage_7_0_t280;
    FSM_dct_8x8_stage_7_0_t282 = FSM_dct_8x8_stage_7_0_t281[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t283 = FSM_dct_8x8_stage_7_0_t273;
    FSM_dct_8x8_stage_7_0_t283[FSM_dct_8x8_stage_7_0_t276 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t282;
    FSM_dct_8x8_stage_7_0_t284 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_7_0_t285 = FSM_dct_8x8_stage_7_0_t284[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t286 = FSM_dct_8x8_stage_7_0_t285[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t287 = FSM_dct_8x8_stage_7_0_t283;
    FSM_dct_8x8_stage_7_0_t287[FSM_dct_8x8_stage_7_0_t286 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t280;
    FSM_dct_8x8_stage_7_0_t288 = 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_7_0_t289 = FSM_dct_8x8_stage_7_0_t288[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t290 = 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_7_0_t291 = FSM_dct_8x8_stage_7_0_t290[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t292 = i_data_in[FSM_dct_8x8_stage_7_0_t291 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t293 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_7_0_t294 = FSM_dct_8x8_stage_7_0_t293[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t295 = FSM_dct_8x8_stage_7_0_t294[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t296 = i_data_in[FSM_dct_8x8_stage_7_0_t295 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t297 = FSM_dct_8x8_stage_7_0_t292 + FSM_dct_8x8_stage_7_0_t296;
    FSM_dct_8x8_stage_7_0_t298 = FSM_dct_8x8_stage_7_0_t297[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t299 = FSM_dct_8x8_stage_7_0_t287;
    FSM_dct_8x8_stage_7_0_t299[FSM_dct_8x8_stage_7_0_t289 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t298;
    FSM_dct_8x8_stage_7_0_t300 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_7_0_t301 = FSM_dct_8x8_stage_7_0_t300[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t302 = FSM_dct_8x8_stage_7_0_t301[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t303 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_7_0_t304 = FSM_dct_8x8_stage_7_0_t303[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t305 = FSM_dct_8x8_stage_7_0_t304[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t306 = i_data_in[FSM_dct_8x8_stage_7_0_t305 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t307 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_7_0_t308 = FSM_dct_8x8_stage_7_0_t307[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t309 = FSM_dct_8x8_stage_7_0_t308[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t310 = i_data_in[FSM_dct_8x8_stage_7_0_t309 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t311 = FSM_dct_8x8_stage_7_0_t306 + FSM_dct_8x8_stage_7_0_t310;
    FSM_dct_8x8_stage_7_0_t312 = FSM_dct_8x8_stage_7_0_t311[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t313 = FSM_dct_8x8_stage_7_0_t299;
    FSM_dct_8x8_stage_7_0_t313[FSM_dct_8x8_stage_7_0_t302 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t312;
    FSM_dct_8x8_stage_7_0_t314 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_7_0_t315 = FSM_dct_8x8_stage_7_0_t314[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t316 = FSM_dct_8x8_stage_7_0_t315[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t317 = FSM_dct_8x8_stage_7_0_t313;
    FSM_dct_8x8_stage_7_0_t317[FSM_dct_8x8_stage_7_0_t316 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t306 - FSM_dct_8x8_stage_7_0_t310;
    FSM_dct_8x8_stage_7_0_t318 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_7_0_t319 = FSM_dct_8x8_stage_7_0_t318[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t320 = FSM_dct_8x8_stage_7_0_t319[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t321 = FSM_dct_8x8_stage_7_0_t317;
    FSM_dct_8x8_stage_7_0_t321[FSM_dct_8x8_stage_7_0_t320 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t292 - FSM_dct_8x8_stage_7_0_t296;
    FSM_dct_8x8_stage_7_0_t322 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_7_0_t323 = FSM_dct_8x8_stage_7_0_t322[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t324 = FSM_dct_8x8_stage_7_0_t323[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t325 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_7_0_t326 = FSM_dct_8x8_stage_7_0_t325[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t327 = FSM_dct_8x8_stage_7_0_t326[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t328 = i_data_in[FSM_dct_8x8_stage_7_0_t327 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t329 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_7_0_t330 = FSM_dct_8x8_stage_7_0_t329[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t331 = FSM_dct_8x8_stage_7_0_t330[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t332 = i_data_in[FSM_dct_8x8_stage_7_0_t331 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t333 = FSM_dct_8x8_stage_7_0_t328 + FSM_dct_8x8_stage_7_0_t332;
    FSM_dct_8x8_stage_7_0_t334 = FSM_dct_8x8_stage_7_0_t333[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t335 = FSM_dct_8x8_stage_7_0_t321;
    FSM_dct_8x8_stage_7_0_t335[FSM_dct_8x8_stage_7_0_t324 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t334;
    FSM_dct_8x8_stage_7_0_t336 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_7_0_t337 = FSM_dct_8x8_stage_7_0_t336[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t338 = FSM_dct_8x8_stage_7_0_t337[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t339 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_7_0_t340 = FSM_dct_8x8_stage_7_0_t339[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t341 = FSM_dct_8x8_stage_7_0_t340[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t342 = i_data_in[FSM_dct_8x8_stage_7_0_t341 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t343 = FSM_dct_8x8_stage_7_0_t332 + FSM_dct_8x8_stage_7_0_t342;
    FSM_dct_8x8_stage_7_0_t344 = FSM_dct_8x8_stage_7_0_t343[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t345 = FSM_dct_8x8_stage_7_0_t335;
    FSM_dct_8x8_stage_7_0_t345[FSM_dct_8x8_stage_7_0_t338 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t344;
    FSM_dct_8x8_stage_7_0_t346 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_7_0_t347 = FSM_dct_8x8_stage_7_0_t346[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t348 = FSM_dct_8x8_stage_7_0_t347[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t349 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_7_0_t350 = FSM_dct_8x8_stage_7_0_t349[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t351 = FSM_dct_8x8_stage_7_0_t350[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t352 = i_data_in[FSM_dct_8x8_stage_7_0_t351 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t353 = FSM_dct_8x8_stage_7_0_t342 + FSM_dct_8x8_stage_7_0_t352;
    FSM_dct_8x8_stage_7_0_t354 = FSM_dct_8x8_stage_7_0_t353[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t355 = FSM_dct_8x8_stage_7_0_t345;
    FSM_dct_8x8_stage_7_0_t355[FSM_dct_8x8_stage_7_0_t348 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t354;
    FSM_dct_8x8_stage_7_0_t356 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_7_0_t357 = FSM_dct_8x8_stage_7_0_t356[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t358 = FSM_dct_8x8_stage_7_0_t357[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t359 = FSM_dct_8x8_stage_7_0_t355;
    FSM_dct_8x8_stage_7_0_t359[FSM_dct_8x8_stage_7_0_t358 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t352;
    FSM_dct_8x8_stage_7_0_t360 = 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_7_0_t361 = FSM_dct_8x8_stage_7_0_t360[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t362 = 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_7_0_t363 = FSM_dct_8x8_stage_7_0_t362[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t364 = i_data_in[FSM_dct_8x8_stage_7_0_t363 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t365 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_7_0_t366 = FSM_dct_8x8_stage_7_0_t365[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t367 = FSM_dct_8x8_stage_7_0_t366[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t368 = i_data_in[FSM_dct_8x8_stage_7_0_t367 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t369 = FSM_dct_8x8_stage_7_0_t364 + FSM_dct_8x8_stage_7_0_t368;
    FSM_dct_8x8_stage_7_0_t370 = FSM_dct_8x8_stage_7_0_t369[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t371 = FSM_dct_8x8_stage_7_0_t359;
    FSM_dct_8x8_stage_7_0_t371[FSM_dct_8x8_stage_7_0_t361 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t370;
    FSM_dct_8x8_stage_7_0_t372 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_7_0_t373 = FSM_dct_8x8_stage_7_0_t372[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t374 = FSM_dct_8x8_stage_7_0_t373[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t375 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_7_0_t376 = FSM_dct_8x8_stage_7_0_t375[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t377 = FSM_dct_8x8_stage_7_0_t376[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t378 = i_data_in[FSM_dct_8x8_stage_7_0_t377 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t379 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_7_0_t380 = FSM_dct_8x8_stage_7_0_t379[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t381 = FSM_dct_8x8_stage_7_0_t380[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t382 = i_data_in[FSM_dct_8x8_stage_7_0_t381 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t383 = FSM_dct_8x8_stage_7_0_t378 + FSM_dct_8x8_stage_7_0_t382;
    FSM_dct_8x8_stage_7_0_t384 = FSM_dct_8x8_stage_7_0_t383[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t385 = FSM_dct_8x8_stage_7_0_t371;
    FSM_dct_8x8_stage_7_0_t385[FSM_dct_8x8_stage_7_0_t374 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t384;
    FSM_dct_8x8_stage_7_0_t386 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_7_0_t387 = FSM_dct_8x8_stage_7_0_t386[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t388 = FSM_dct_8x8_stage_7_0_t387[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t389 = FSM_dct_8x8_stage_7_0_t385;
    FSM_dct_8x8_stage_7_0_t389[FSM_dct_8x8_stage_7_0_t388 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t378 - FSM_dct_8x8_stage_7_0_t382;
    FSM_dct_8x8_stage_7_0_t390 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_7_0_t391 = FSM_dct_8x8_stage_7_0_t390[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t392 = FSM_dct_8x8_stage_7_0_t391[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t393 = FSM_dct_8x8_stage_7_0_t389;
    FSM_dct_8x8_stage_7_0_t393[FSM_dct_8x8_stage_7_0_t392 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t364 - FSM_dct_8x8_stage_7_0_t368;
    FSM_dct_8x8_stage_7_0_t394 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_7_0_t395 = FSM_dct_8x8_stage_7_0_t394[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t396 = FSM_dct_8x8_stage_7_0_t395[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t397 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_7_0_t398 = FSM_dct_8x8_stage_7_0_t397[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t399 = FSM_dct_8x8_stage_7_0_t398[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t400 = i_data_in[FSM_dct_8x8_stage_7_0_t399 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t401 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_7_0_t402 = FSM_dct_8x8_stage_7_0_t401[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t403 = FSM_dct_8x8_stage_7_0_t402[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t404 = i_data_in[FSM_dct_8x8_stage_7_0_t403 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t405 = FSM_dct_8x8_stage_7_0_t400 + FSM_dct_8x8_stage_7_0_t404;
    FSM_dct_8x8_stage_7_0_t406 = FSM_dct_8x8_stage_7_0_t405[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t407 = FSM_dct_8x8_stage_7_0_t393;
    FSM_dct_8x8_stage_7_0_t407[FSM_dct_8x8_stage_7_0_t396 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t406;
    FSM_dct_8x8_stage_7_0_t408 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_7_0_t409 = FSM_dct_8x8_stage_7_0_t408[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t410 = FSM_dct_8x8_stage_7_0_t409[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t411 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_7_0_t412 = FSM_dct_8x8_stage_7_0_t411[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t413 = FSM_dct_8x8_stage_7_0_t412[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t414 = i_data_in[FSM_dct_8x8_stage_7_0_t413 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t415 = FSM_dct_8x8_stage_7_0_t404 + FSM_dct_8x8_stage_7_0_t414;
    FSM_dct_8x8_stage_7_0_t416 = FSM_dct_8x8_stage_7_0_t415[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t417 = FSM_dct_8x8_stage_7_0_t407;
    FSM_dct_8x8_stage_7_0_t417[FSM_dct_8x8_stage_7_0_t410 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t416;
    FSM_dct_8x8_stage_7_0_t418 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_7_0_t419 = FSM_dct_8x8_stage_7_0_t418[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t420 = FSM_dct_8x8_stage_7_0_t419[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t421 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_7_0_t422 = FSM_dct_8x8_stage_7_0_t421[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t423 = FSM_dct_8x8_stage_7_0_t422[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t424 = i_data_in[FSM_dct_8x8_stage_7_0_t423 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t425 = FSM_dct_8x8_stage_7_0_t414 + FSM_dct_8x8_stage_7_0_t424;
    FSM_dct_8x8_stage_7_0_t426 = FSM_dct_8x8_stage_7_0_t425[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t427 = FSM_dct_8x8_stage_7_0_t417;
    FSM_dct_8x8_stage_7_0_t427[FSM_dct_8x8_stage_7_0_t420 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t426;
    FSM_dct_8x8_stage_7_0_t428 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_7_0_t429 = FSM_dct_8x8_stage_7_0_t428[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t430 = FSM_dct_8x8_stage_7_0_t429[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t431 = FSM_dct_8x8_stage_7_0_t427;
    FSM_dct_8x8_stage_7_0_t431[FSM_dct_8x8_stage_7_0_t430 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t424;
    FSM_dct_8x8_stage_7_0_t432 = 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_7_0_t433 = FSM_dct_8x8_stage_7_0_t432[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t434 = 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_7_0_t435 = FSM_dct_8x8_stage_7_0_t434[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t436 = i_data_in[FSM_dct_8x8_stage_7_0_t435 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t437 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_7_0_t438 = FSM_dct_8x8_stage_7_0_t437[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t439 = FSM_dct_8x8_stage_7_0_t438[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t440 = i_data_in[FSM_dct_8x8_stage_7_0_t439 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t441 = FSM_dct_8x8_stage_7_0_t436 + FSM_dct_8x8_stage_7_0_t440;
    FSM_dct_8x8_stage_7_0_t442 = FSM_dct_8x8_stage_7_0_t441[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t443 = FSM_dct_8x8_stage_7_0_t431;
    FSM_dct_8x8_stage_7_0_t443[FSM_dct_8x8_stage_7_0_t433 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t442;
    FSM_dct_8x8_stage_7_0_t444 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_7_0_t445 = FSM_dct_8x8_stage_7_0_t444[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t446 = FSM_dct_8x8_stage_7_0_t445[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t447 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_7_0_t448 = FSM_dct_8x8_stage_7_0_t447[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t449 = FSM_dct_8x8_stage_7_0_t448[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t450 = i_data_in[FSM_dct_8x8_stage_7_0_t449 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t451 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_7_0_t452 = FSM_dct_8x8_stage_7_0_t451[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t453 = FSM_dct_8x8_stage_7_0_t452[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t454 = i_data_in[FSM_dct_8x8_stage_7_0_t453 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t455 = FSM_dct_8x8_stage_7_0_t450 + FSM_dct_8x8_stage_7_0_t454;
    FSM_dct_8x8_stage_7_0_t456 = FSM_dct_8x8_stage_7_0_t455[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t457 = FSM_dct_8x8_stage_7_0_t443;
    FSM_dct_8x8_stage_7_0_t457[FSM_dct_8x8_stage_7_0_t446 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t456;
    FSM_dct_8x8_stage_7_0_t458 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_7_0_t459 = FSM_dct_8x8_stage_7_0_t458[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t460 = FSM_dct_8x8_stage_7_0_t459[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t461 = FSM_dct_8x8_stage_7_0_t457;
    FSM_dct_8x8_stage_7_0_t461[FSM_dct_8x8_stage_7_0_t460 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t450 - FSM_dct_8x8_stage_7_0_t454;
    FSM_dct_8x8_stage_7_0_t462 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_7_0_t463 = FSM_dct_8x8_stage_7_0_t462[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t464 = FSM_dct_8x8_stage_7_0_t463[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t465 = FSM_dct_8x8_stage_7_0_t461;
    FSM_dct_8x8_stage_7_0_t465[FSM_dct_8x8_stage_7_0_t464 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t436 - FSM_dct_8x8_stage_7_0_t440;
    FSM_dct_8x8_stage_7_0_t466 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_7_0_t467 = FSM_dct_8x8_stage_7_0_t466[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t468 = FSM_dct_8x8_stage_7_0_t467[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t469 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_7_0_t470 = FSM_dct_8x8_stage_7_0_t469[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t471 = FSM_dct_8x8_stage_7_0_t470[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t472 = i_data_in[FSM_dct_8x8_stage_7_0_t471 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t473 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_7_0_t474 = FSM_dct_8x8_stage_7_0_t473[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t475 = FSM_dct_8x8_stage_7_0_t474[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t476 = i_data_in[FSM_dct_8x8_stage_7_0_t475 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t477 = FSM_dct_8x8_stage_7_0_t472 + FSM_dct_8x8_stage_7_0_t476;
    FSM_dct_8x8_stage_7_0_t478 = FSM_dct_8x8_stage_7_0_t477[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t479 = FSM_dct_8x8_stage_7_0_t465;
    FSM_dct_8x8_stage_7_0_t479[FSM_dct_8x8_stage_7_0_t468 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t478;
    FSM_dct_8x8_stage_7_0_t480 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_7_0_t481 = FSM_dct_8x8_stage_7_0_t480[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t482 = FSM_dct_8x8_stage_7_0_t481[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t483 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_7_0_t484 = FSM_dct_8x8_stage_7_0_t483[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t485 = FSM_dct_8x8_stage_7_0_t484[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t486 = i_data_in[FSM_dct_8x8_stage_7_0_t485 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t487 = FSM_dct_8x8_stage_7_0_t476 + FSM_dct_8x8_stage_7_0_t486;
    FSM_dct_8x8_stage_7_0_t488 = FSM_dct_8x8_stage_7_0_t487[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t489 = FSM_dct_8x8_stage_7_0_t479;
    FSM_dct_8x8_stage_7_0_t489[FSM_dct_8x8_stage_7_0_t482 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t488;
    FSM_dct_8x8_stage_7_0_t490 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_7_0_t491 = FSM_dct_8x8_stage_7_0_t490[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t492 = FSM_dct_8x8_stage_7_0_t491[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t493 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_7_0_t494 = FSM_dct_8x8_stage_7_0_t493[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t495 = FSM_dct_8x8_stage_7_0_t494[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t496 = i_data_in[FSM_dct_8x8_stage_7_0_t495 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t497 = FSM_dct_8x8_stage_7_0_t486 + FSM_dct_8x8_stage_7_0_t496;
    FSM_dct_8x8_stage_7_0_t498 = FSM_dct_8x8_stage_7_0_t497[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t499 = FSM_dct_8x8_stage_7_0_t489;
    FSM_dct_8x8_stage_7_0_t499[FSM_dct_8x8_stage_7_0_t492 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t498;
    FSM_dct_8x8_stage_7_0_t500 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_7_0_t501 = FSM_dct_8x8_stage_7_0_t500[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t502 = FSM_dct_8x8_stage_7_0_t501[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t503 = FSM_dct_8x8_stage_7_0_t499;
    FSM_dct_8x8_stage_7_0_t503[FSM_dct_8x8_stage_7_0_t502 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t496;
    FSM_dct_8x8_stage_7_0_t504 = 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_7_0_t505 = FSM_dct_8x8_stage_7_0_t504[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t506 = 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_7_0_t507 = FSM_dct_8x8_stage_7_0_t506[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t508 = i_data_in[FSM_dct_8x8_stage_7_0_t507 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t509 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_7_0_t510 = FSM_dct_8x8_stage_7_0_t509[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t511 = FSM_dct_8x8_stage_7_0_t510[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t512 = i_data_in[FSM_dct_8x8_stage_7_0_t511 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t513 = FSM_dct_8x8_stage_7_0_t508 + FSM_dct_8x8_stage_7_0_t512;
    FSM_dct_8x8_stage_7_0_t514 = FSM_dct_8x8_stage_7_0_t513[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t515 = FSM_dct_8x8_stage_7_0_t503;
    FSM_dct_8x8_stage_7_0_t515[FSM_dct_8x8_stage_7_0_t505 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t514;
    FSM_dct_8x8_stage_7_0_t516 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_7_0_t517 = FSM_dct_8x8_stage_7_0_t516[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t518 = FSM_dct_8x8_stage_7_0_t517[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t519 = 32'b00000000000000000000000000001000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_7_0_t520 = FSM_dct_8x8_stage_7_0_t519[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t521 = FSM_dct_8x8_stage_7_0_t520[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t522 = i_data_in[FSM_dct_8x8_stage_7_0_t521 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t523 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_7_0_t524 = FSM_dct_8x8_stage_7_0_t523[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t525 = FSM_dct_8x8_stage_7_0_t524[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t526 = i_data_in[FSM_dct_8x8_stage_7_0_t525 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t527 = FSM_dct_8x8_stage_7_0_t522 + FSM_dct_8x8_stage_7_0_t526;
    FSM_dct_8x8_stage_7_0_t528 = FSM_dct_8x8_stage_7_0_t527[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t529 = FSM_dct_8x8_stage_7_0_t515;
    FSM_dct_8x8_stage_7_0_t529[FSM_dct_8x8_stage_7_0_t518 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t528;
    FSM_dct_8x8_stage_7_0_t530 = 32'b00000000000000000000000000010000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_7_0_t531 = FSM_dct_8x8_stage_7_0_t530[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t532 = FSM_dct_8x8_stage_7_0_t531[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t533 = FSM_dct_8x8_stage_7_0_t529;
    FSM_dct_8x8_stage_7_0_t533[FSM_dct_8x8_stage_7_0_t532 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t522 - FSM_dct_8x8_stage_7_0_t526;
    FSM_dct_8x8_stage_7_0_t534 = 32'b00000000000000000000000000011000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_7_0_t535 = FSM_dct_8x8_stage_7_0_t534[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t536 = FSM_dct_8x8_stage_7_0_t535[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t537 = FSM_dct_8x8_stage_7_0_t533;
    FSM_dct_8x8_stage_7_0_t537[FSM_dct_8x8_stage_7_0_t536 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t508 - FSM_dct_8x8_stage_7_0_t512;
    FSM_dct_8x8_stage_7_0_t538 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_7_0_t539 = FSM_dct_8x8_stage_7_0_t538[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t540 = FSM_dct_8x8_stage_7_0_t539[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t541 = 32'b00000000000000000000000000100000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_7_0_t542 = FSM_dct_8x8_stage_7_0_t541[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t543 = FSM_dct_8x8_stage_7_0_t542[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t544 = i_data_in[FSM_dct_8x8_stage_7_0_t543 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t545 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_7_0_t546 = FSM_dct_8x8_stage_7_0_t545[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t547 = FSM_dct_8x8_stage_7_0_t546[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t548 = i_data_in[FSM_dct_8x8_stage_7_0_t547 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t549 = FSM_dct_8x8_stage_7_0_t544 + FSM_dct_8x8_stage_7_0_t548;
    FSM_dct_8x8_stage_7_0_t550 = FSM_dct_8x8_stage_7_0_t549[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t551 = FSM_dct_8x8_stage_7_0_t537;
    FSM_dct_8x8_stage_7_0_t551[FSM_dct_8x8_stage_7_0_t540 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t550;
    FSM_dct_8x8_stage_7_0_t552 = 32'b00000000000000000000000000101000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_7_0_t553 = FSM_dct_8x8_stage_7_0_t552[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t554 = FSM_dct_8x8_stage_7_0_t553[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t555 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_7_0_t556 = FSM_dct_8x8_stage_7_0_t555[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t557 = FSM_dct_8x8_stage_7_0_t556[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t558 = i_data_in[FSM_dct_8x8_stage_7_0_t557 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t559 = FSM_dct_8x8_stage_7_0_t548 + FSM_dct_8x8_stage_7_0_t558;
    FSM_dct_8x8_stage_7_0_t560 = FSM_dct_8x8_stage_7_0_t559[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t561 = FSM_dct_8x8_stage_7_0_t551;
    FSM_dct_8x8_stage_7_0_t561[FSM_dct_8x8_stage_7_0_t554 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t560;
    FSM_dct_8x8_stage_7_0_t562 = 32'b00000000000000000000000000110000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_7_0_t563 = FSM_dct_8x8_stage_7_0_t562[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t564 = FSM_dct_8x8_stage_7_0_t563[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t565 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_7_0_t566 = FSM_dct_8x8_stage_7_0_t565[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t567 = FSM_dct_8x8_stage_7_0_t566[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t568 = i_data_in[FSM_dct_8x8_stage_7_0_t567 * 32 +: 32];
    FSM_dct_8x8_stage_7_0_t569 = FSM_dct_8x8_stage_7_0_t558 + FSM_dct_8x8_stage_7_0_t568;
    FSM_dct_8x8_stage_7_0_t570 = FSM_dct_8x8_stage_7_0_t569[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t571 = FSM_dct_8x8_stage_7_0_t561;
    FSM_dct_8x8_stage_7_0_t571[FSM_dct_8x8_stage_7_0_t564 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t570;
    FSM_dct_8x8_stage_7_0_t572 = 32'b00000000000000000000000000111000 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_7_0_t573 = FSM_dct_8x8_stage_7_0_t572[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_7_0_t574 = FSM_dct_8x8_stage_7_0_t573[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_7_0_t575 = FSM_dct_8x8_stage_7_0_t571;
    FSM_dct_8x8_stage_7_0_t575[FSM_dct_8x8_stage_7_0_t574 * 32 +: 32] = FSM_dct_8x8_stage_7_0_t568;
end

assign FSM_dct_8x8_stage_7_0_in_ready = 1'b1;

always @(posedge clk) begin
    FSM_dct_8x8_stage_7_0_st_dummy_reg <= FSM_dct_8x8_stage_7_0_st_dummy_reg;
    if (rst) begin
        FSM_dct_8x8_stage_7_0_st_dummy_reg <= 32'b0;
    end
end
/* End submodules of dct_8x8_stage_7 */
/* End module dct_8x8_stage_7 */
endgenerate
endmodule
