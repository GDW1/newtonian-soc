`timescale 1ns / 1ps

module dct_8x8_stage_4_inner
(
    input wire clk,
    input wire rst,
    input wire [2048-1:0] i_data_in,
    input wire i_valid,
    output wire i_ready,
    output wire [2048-1:0] o_data_out,
    output wire o_valid,
    input wire o_ready
);

generate
/*
    Begin module dct_8x8_stage_4
*/
/*
    Wires declared by dct_8x8_stage_4
*/
wire FSM_dct_8x8_stage_4_0_in_ready;
wire FSM_dct_8x8_stage_4_0_out_valid;
/* End wires declared by dct_8x8_stage_4 */

/*
    Submodules of dct_8x8_stage_4
*/
reg [32-1:0] FSM_dct_8x8_stage_4_0_st_dummy_reg = 32'b0;

reg [64-1:0] FSM_dct_8x8_stage_4_0_t0;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t1;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t2;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t3;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t4;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t5;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t6;
reg [2048-1:0] FSM_dct_8x8_stage_4_0_t7;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t8;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t9;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t10;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t11;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t12;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t13;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t14;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t15;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t16;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t17;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t18;
reg [2048-1:0] FSM_dct_8x8_stage_4_0_t19;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t20;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t21;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t22;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t23;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t24;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t25;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t26;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t27;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t28;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t29;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t30;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t31;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t32;
reg [2048-1:0] FSM_dct_8x8_stage_4_0_t33;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t34;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t35;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t36;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t37;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t38;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t39;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t40;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t41;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t42;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t43;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t44;
reg [2048-1:0] FSM_dct_8x8_stage_4_0_t45;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t46;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t47;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t48;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t49;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t50;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t51;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t52;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t53;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t54;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t55;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t56;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t57;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t58;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t59;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t60;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t61;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t62;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t63;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t64;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t65;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t66;
reg [2048-1:0] FSM_dct_8x8_stage_4_0_t67;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t68;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t69;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t70;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t71;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t72;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t73;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t74;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t75;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t76;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t77;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t78;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t79;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t80;
reg [2048-1:0] FSM_dct_8x8_stage_4_0_t81;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t82;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t83;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t84;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t85;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t86;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t87;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t88;
reg [2048-1:0] FSM_dct_8x8_stage_4_0_t89;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t90;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t91;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t92;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t93;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t94;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t95;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t96;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t97;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t98;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t99;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t100;
reg [2048-1:0] FSM_dct_8x8_stage_4_0_t101;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t102;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t103;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t104;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t105;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t106;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t107;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t108;
reg [2048-1:0] FSM_dct_8x8_stage_4_0_t109;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t110;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t111;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t112;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t113;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t114;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t115;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t116;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t117;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t118;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t119;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t120;
reg [2048-1:0] FSM_dct_8x8_stage_4_0_t121;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t122;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t123;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t124;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t125;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t126;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t127;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t128;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t129;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t130;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t131;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t132;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t133;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t134;
reg [2048-1:0] FSM_dct_8x8_stage_4_0_t135;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t136;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t137;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t138;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t139;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t140;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t141;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t142;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t143;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t144;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t145;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t146;
reg [2048-1:0] FSM_dct_8x8_stage_4_0_t147;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t148;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t149;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t150;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t151;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t152;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t153;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t154;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t155;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t156;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t157;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t158;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t159;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t160;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t161;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t162;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t163;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t164;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t165;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t166;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t167;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t168;
reg [2048-1:0] FSM_dct_8x8_stage_4_0_t169;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t170;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t171;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t172;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t173;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t174;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t175;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t176;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t177;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t178;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t179;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t180;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t181;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t182;
reg [2048-1:0] FSM_dct_8x8_stage_4_0_t183;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t184;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t185;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t186;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t187;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t188;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t189;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t190;
reg [2048-1:0] FSM_dct_8x8_stage_4_0_t191;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t192;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t193;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t194;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t195;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t196;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t197;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t198;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t199;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t200;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t201;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t202;
reg [2048-1:0] FSM_dct_8x8_stage_4_0_t203;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t204;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t205;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t206;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t207;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t208;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t209;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t210;
reg [2048-1:0] FSM_dct_8x8_stage_4_0_t211;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t212;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t213;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t214;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t215;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t216;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t217;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t218;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t219;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t220;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t221;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t222;
reg [2048-1:0] FSM_dct_8x8_stage_4_0_t223;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t224;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t225;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t226;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t227;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t228;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t229;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t230;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t231;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t232;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t233;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t234;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t235;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t236;
reg [2048-1:0] FSM_dct_8x8_stage_4_0_t237;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t238;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t239;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t240;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t241;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t242;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t243;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t244;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t245;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t246;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t247;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t248;
reg [2048-1:0] FSM_dct_8x8_stage_4_0_t249;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t250;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t251;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t252;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t253;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t254;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t255;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t256;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t257;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t258;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t259;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t260;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t261;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t262;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t263;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t264;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t265;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t266;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t267;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t268;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t269;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t270;
reg [2048-1:0] FSM_dct_8x8_stage_4_0_t271;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t272;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t273;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t274;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t275;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t276;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t277;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t278;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t279;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t280;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t281;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t282;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t283;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t284;
reg [2048-1:0] FSM_dct_8x8_stage_4_0_t285;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t286;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t287;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t288;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t289;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t290;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t291;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t292;
reg [2048-1:0] FSM_dct_8x8_stage_4_0_t293;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t294;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t295;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t296;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t297;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t298;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t299;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t300;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t301;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t302;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t303;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t304;
reg [2048-1:0] FSM_dct_8x8_stage_4_0_t305;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t306;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t307;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t308;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t309;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t310;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t311;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t312;
reg [2048-1:0] FSM_dct_8x8_stage_4_0_t313;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t314;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t315;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t316;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t317;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t318;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t319;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t320;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t321;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t322;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t323;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t324;
reg [2048-1:0] FSM_dct_8x8_stage_4_0_t325;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t326;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t327;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t328;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t329;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t330;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t331;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t332;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t333;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t334;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t335;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t336;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t337;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t338;
reg [2048-1:0] FSM_dct_8x8_stage_4_0_t339;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t340;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t341;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t342;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t343;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t344;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t345;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t346;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t347;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t348;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t349;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t350;
reg [2048-1:0] FSM_dct_8x8_stage_4_0_t351;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t352;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t353;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t354;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t355;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t356;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t357;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t358;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t359;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t360;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t361;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t362;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t363;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t364;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t365;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t366;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t367;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t368;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t369;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t370;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t371;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t372;
reg [2048-1:0] FSM_dct_8x8_stage_4_0_t373;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t374;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t375;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t376;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t377;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t378;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t379;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t380;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t381;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t382;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t383;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t384;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t385;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t386;
reg [2048-1:0] FSM_dct_8x8_stage_4_0_t387;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t388;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t389;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t390;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t391;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t392;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t393;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t394;
reg [2048-1:0] FSM_dct_8x8_stage_4_0_t395;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t396;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t397;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t398;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t399;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t400;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t401;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t402;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t403;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t404;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t405;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t406;
reg [2048-1:0] FSM_dct_8x8_stage_4_0_t407;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t408;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t409;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t410;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t411;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t412;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t413;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t414;
reg [2048-1:0] FSM_dct_8x8_stage_4_0_t415;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t416;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t417;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t418;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t419;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t420;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t421;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t422;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t423;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t424;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t425;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t426;
reg [2048-1:0] FSM_dct_8x8_stage_4_0_t427;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t428;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t429;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t430;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t431;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t432;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t433;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t434;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t435;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t436;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t437;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t438;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t439;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t440;
reg [2048-1:0] FSM_dct_8x8_stage_4_0_t441;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t442;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t443;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t444;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t445;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t446;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t447;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t448;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t449;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t450;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t451;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t452;
reg [2048-1:0] FSM_dct_8x8_stage_4_0_t453;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t454;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t455;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t456;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t457;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t458;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t459;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t460;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t461;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t462;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t463;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t464;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t465;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t466;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t467;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t468;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t469;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t470;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t471;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t472;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t473;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t474;
reg [2048-1:0] FSM_dct_8x8_stage_4_0_t475;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t476;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t477;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t478;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t479;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t480;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t481;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t482;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t483;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t484;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t485;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t486;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t487;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t488;
reg [2048-1:0] FSM_dct_8x8_stage_4_0_t489;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t490;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t491;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t492;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t493;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t494;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t495;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t496;
reg [2048-1:0] FSM_dct_8x8_stage_4_0_t497;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t498;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t499;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t500;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t501;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t502;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t503;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t504;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t505;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t506;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t507;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t508;
reg [2048-1:0] FSM_dct_8x8_stage_4_0_t509;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t510;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t511;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t512;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t513;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t514;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t515;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t516;
reg [2048-1:0] FSM_dct_8x8_stage_4_0_t517;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t518;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t519;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t520;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t521;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t522;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t523;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t524;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t525;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t526;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t527;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t528;
reg [2048-1:0] FSM_dct_8x8_stage_4_0_t529;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t530;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t531;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t532;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t533;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t534;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t535;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t536;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t537;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t538;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t539;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t540;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t541;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t542;
reg [2048-1:0] FSM_dct_8x8_stage_4_0_t543;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t544;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t545;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t546;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t547;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t548;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t549;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t550;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t551;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t552;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t553;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t554;
reg [2048-1:0] FSM_dct_8x8_stage_4_0_t555;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t556;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t557;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t558;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t559;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t560;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t561;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t562;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t563;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t564;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t565;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t566;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t567;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t568;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t569;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t570;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t571;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t572;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t573;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t574;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t575;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t576;
reg [2048-1:0] FSM_dct_8x8_stage_4_0_t577;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t578;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t579;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t580;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t581;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t582;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t583;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t584;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t585;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t586;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t587;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t588;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t589;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t590;
reg [2048-1:0] FSM_dct_8x8_stage_4_0_t591;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t592;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t593;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t594;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t595;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t596;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t597;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t598;
reg [2048-1:0] FSM_dct_8x8_stage_4_0_t599;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t600;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t601;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t602;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t603;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t604;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t605;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t606;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t607;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t608;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t609;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t610;
reg [2048-1:0] FSM_dct_8x8_stage_4_0_t611;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t612;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t613;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t614;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t615;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t616;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t617;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t618;
reg [2048-1:0] FSM_dct_8x8_stage_4_0_t619;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t620;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t621;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t622;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t623;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t624;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t625;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t626;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t627;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t628;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t629;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t630;
reg [2048-1:0] FSM_dct_8x8_stage_4_0_t631;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t632;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t633;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t634;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t635;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t636;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t637;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t638;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t639;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t640;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t641;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t642;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t643;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t644;
reg [2048-1:0] FSM_dct_8x8_stage_4_0_t645;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t646;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t647;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t648;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t649;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t650;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t651;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t652;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t653;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t654;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t655;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t656;
reg [2048-1:0] FSM_dct_8x8_stage_4_0_t657;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t658;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t659;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t660;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t661;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t662;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t663;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t664;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t665;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t666;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t667;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t668;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t669;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t670;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t671;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t672;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t673;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t674;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t675;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t676;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t677;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t678;
reg [2048-1:0] FSM_dct_8x8_stage_4_0_t679;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t680;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t681;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t682;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t683;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t684;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t685;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t686;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t687;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t688;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t689;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t690;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t691;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t692;
reg [2048-1:0] FSM_dct_8x8_stage_4_0_t693;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t694;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t695;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t696;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t697;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t698;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t699;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t700;
reg [2048-1:0] FSM_dct_8x8_stage_4_0_t701;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t702;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t703;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t704;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t705;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t706;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t707;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t708;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t709;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t710;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t711;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t712;
reg [2048-1:0] FSM_dct_8x8_stage_4_0_t713;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t714;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t715;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t716;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t717;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t718;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t719;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t720;
reg [2048-1:0] FSM_dct_8x8_stage_4_0_t721;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t722;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t723;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t724;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t725;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t726;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t727;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t728;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t729;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t730;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t731;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t732;
reg [2048-1:0] FSM_dct_8x8_stage_4_0_t733;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t734;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t735;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t736;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t737;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t738;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t739;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t740;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t741;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t742;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t743;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t744;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t745;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t746;
reg [2048-1:0] FSM_dct_8x8_stage_4_0_t747;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t748;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t749;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t750;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t751;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t752;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t753;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t754;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t755;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t756;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t757;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t758;
reg [2048-1:0] FSM_dct_8x8_stage_4_0_t759;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t760;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t761;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t762;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t763;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t764;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t765;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t766;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t767;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t768;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t769;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t770;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t771;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t772;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t773;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t774;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t775;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t776;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t777;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t778;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t779;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t780;
reg [2048-1:0] FSM_dct_8x8_stage_4_0_t781;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t782;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t783;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t784;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t785;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t786;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t787;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t788;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t789;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t790;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t791;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t792;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t793;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t794;
reg [2048-1:0] FSM_dct_8x8_stage_4_0_t795;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t796;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t797;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t798;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t799;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t800;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t801;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t802;
reg [2048-1:0] FSM_dct_8x8_stage_4_0_t803;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t804;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t805;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t806;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t807;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t808;
reg [64-1:0] FSM_dct_8x8_stage_4_0_t809;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t810;
reg [33-1:0] FSM_dct_8x8_stage_4_0_t811;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t812;
reg [6-1:0] FSM_dct_8x8_stage_4_0_t813;
reg [32-1:0] FSM_dct_8x8_stage_4_0_t814;
reg [2048-1:0] FSM_dct_8x8_stage_4_0_t815;

/*
    Wiring by dct_8x8_stage_4
*/
assign i_ready = FSM_dct_8x8_stage_4_0_in_ready;
assign o_data_out = FSM_dct_8x8_stage_4_0_t815;
assign o_valid = FSM_dct_8x8_stage_4_0_out_valid;
/* End wiring by dct_8x8_stage_4 */

assign FSM_dct_8x8_stage_4_0_out_valid = 1'b1;

initial begin
    FSM_dct_8x8_stage_4_0_t0 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_4_0_t1 = FSM_dct_8x8_stage_4_0_t0[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t2 = FSM_dct_8x8_stage_4_0_t1[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t3 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_4_0_t4 = FSM_dct_8x8_stage_4_0_t3[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t5 = FSM_dct_8x8_stage_4_0_t4[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t6 = i_data_in[FSM_dct_8x8_stage_4_0_t5 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t7 = 2048'b0;
    FSM_dct_8x8_stage_4_0_t7[FSM_dct_8x8_stage_4_0_t2 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t6;
    FSM_dct_8x8_stage_4_0_t8 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_4_0_t9 = FSM_dct_8x8_stage_4_0_t8[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t10 = FSM_dct_8x8_stage_4_0_t9 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_4_0_t11 = FSM_dct_8x8_stage_4_0_t10[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t12 = FSM_dct_8x8_stage_4_0_t11[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t13 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_4_0_t14 = FSM_dct_8x8_stage_4_0_t13[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t15 = FSM_dct_8x8_stage_4_0_t14 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_4_0_t16 = FSM_dct_8x8_stage_4_0_t15[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t17 = FSM_dct_8x8_stage_4_0_t16[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t18 = i_data_in[FSM_dct_8x8_stage_4_0_t17 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t19 = FSM_dct_8x8_stage_4_0_t7;
    FSM_dct_8x8_stage_4_0_t19[FSM_dct_8x8_stage_4_0_t12 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t18;
    FSM_dct_8x8_stage_4_0_t20 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_4_0_t21 = FSM_dct_8x8_stage_4_0_t20[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t22 = FSM_dct_8x8_stage_4_0_t21 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_4_0_t23 = FSM_dct_8x8_stage_4_0_t22[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t24 = FSM_dct_8x8_stage_4_0_t23[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t25 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_4_0_t26 = FSM_dct_8x8_stage_4_0_t25[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t27 = FSM_dct_8x8_stage_4_0_t26 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_4_0_t28 = FSM_dct_8x8_stage_4_0_t27[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t29 = FSM_dct_8x8_stage_4_0_t28[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t30 = i_data_in[FSM_dct_8x8_stage_4_0_t29 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t31 = FSM_dct_8x8_stage_4_0_t30 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t32 = FSM_dct_8x8_stage_4_0_t31[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t33 = FSM_dct_8x8_stage_4_0_t19;
    FSM_dct_8x8_stage_4_0_t33[FSM_dct_8x8_stage_4_0_t24 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t32;
    FSM_dct_8x8_stage_4_0_t34 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_4_0_t35 = FSM_dct_8x8_stage_4_0_t34[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t36 = FSM_dct_8x8_stage_4_0_t35 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_4_0_t37 = FSM_dct_8x8_stage_4_0_t36[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t38 = FSM_dct_8x8_stage_4_0_t37[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t39 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_4_0_t40 = FSM_dct_8x8_stage_4_0_t39[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t41 = FSM_dct_8x8_stage_4_0_t40 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_4_0_t42 = FSM_dct_8x8_stage_4_0_t41[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t43 = FSM_dct_8x8_stage_4_0_t42[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t44 = i_data_in[FSM_dct_8x8_stage_4_0_t43 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t45 = FSM_dct_8x8_stage_4_0_t33;
    FSM_dct_8x8_stage_4_0_t45[FSM_dct_8x8_stage_4_0_t38 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t44;
    FSM_dct_8x8_stage_4_0_t46 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_4_0_t47 = FSM_dct_8x8_stage_4_0_t46[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t48 = FSM_dct_8x8_stage_4_0_t47 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_4_0_t49 = FSM_dct_8x8_stage_4_0_t48[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t50 = FSM_dct_8x8_stage_4_0_t49[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t51 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_4_0_t52 = FSM_dct_8x8_stage_4_0_t51[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t53 = FSM_dct_8x8_stage_4_0_t52 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_4_0_t54 = FSM_dct_8x8_stage_4_0_t53[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t55 = FSM_dct_8x8_stage_4_0_t54[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t56 = i_data_in[FSM_dct_8x8_stage_4_0_t55 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t57 = FSM_dct_8x8_stage_4_0_t56 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t58 = FSM_dct_8x8_stage_4_0_t57[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t59 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_4_0_t60 = FSM_dct_8x8_stage_4_0_t59[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t61 = FSM_dct_8x8_stage_4_0_t60 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_4_0_t62 = FSM_dct_8x8_stage_4_0_t61[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t63 = FSM_dct_8x8_stage_4_0_t62[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t64 = i_data_in[FSM_dct_8x8_stage_4_0_t63 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t65 = (FSM_dct_8x8_stage_4_0_t64 - FSM_dct_8x8_stage_4_0_t56) * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t66 = FSM_dct_8x8_stage_4_0_t65[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t67 = FSM_dct_8x8_stage_4_0_t45;
    FSM_dct_8x8_stage_4_0_t67[FSM_dct_8x8_stage_4_0_t50 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t58 - FSM_dct_8x8_stage_4_0_t66;
    FSM_dct_8x8_stage_4_0_t68 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_4_0_t69 = FSM_dct_8x8_stage_4_0_t68[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t70 = FSM_dct_8x8_stage_4_0_t69 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_4_0_t71 = FSM_dct_8x8_stage_4_0_t70[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t72 = FSM_dct_8x8_stage_4_0_t71[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t73 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_4_0_t74 = FSM_dct_8x8_stage_4_0_t73[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t75 = FSM_dct_8x8_stage_4_0_t74 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_4_0_t76 = FSM_dct_8x8_stage_4_0_t75[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t77 = FSM_dct_8x8_stage_4_0_t76[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t78 = i_data_in[FSM_dct_8x8_stage_4_0_t77 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t79 = FSM_dct_8x8_stage_4_0_t78 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t80 = FSM_dct_8x8_stage_4_0_t79[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t81 = FSM_dct_8x8_stage_4_0_t67;
    FSM_dct_8x8_stage_4_0_t81[FSM_dct_8x8_stage_4_0_t72 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t80;
    FSM_dct_8x8_stage_4_0_t82 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_4_0_t83 = FSM_dct_8x8_stage_4_0_t82[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t84 = FSM_dct_8x8_stage_4_0_t83 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_4_0_t85 = FSM_dct_8x8_stage_4_0_t84[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t86 = FSM_dct_8x8_stage_4_0_t85[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t87 = FSM_dct_8x8_stage_4_0_t64 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t88 = FSM_dct_8x8_stage_4_0_t87[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t89 = FSM_dct_8x8_stage_4_0_t81;
    FSM_dct_8x8_stage_4_0_t89[FSM_dct_8x8_stage_4_0_t86 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t88 - FSM_dct_8x8_stage_4_0_t66;
    FSM_dct_8x8_stage_4_0_t90 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_4_0_t91 = FSM_dct_8x8_stage_4_0_t90[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t92 = FSM_dct_8x8_stage_4_0_t91 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_4_0_t93 = FSM_dct_8x8_stage_4_0_t92[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t94 = FSM_dct_8x8_stage_4_0_t93[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t95 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_4_0_t96 = FSM_dct_8x8_stage_4_0_t95[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t97 = FSM_dct_8x8_stage_4_0_t96 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_4_0_t98 = FSM_dct_8x8_stage_4_0_t97[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t99 = FSM_dct_8x8_stage_4_0_t98[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t100 = i_data_in[FSM_dct_8x8_stage_4_0_t99 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t101 = FSM_dct_8x8_stage_4_0_t89;
    FSM_dct_8x8_stage_4_0_t101[FSM_dct_8x8_stage_4_0_t94 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t100;
    FSM_dct_8x8_stage_4_0_t102 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_4_0_t103 = FSM_dct_8x8_stage_4_0_t102[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t104 = FSM_dct_8x8_stage_4_0_t103[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t105 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_4_0_t106 = FSM_dct_8x8_stage_4_0_t105[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t107 = FSM_dct_8x8_stage_4_0_t106[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t108 = i_data_in[FSM_dct_8x8_stage_4_0_t107 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t109 = FSM_dct_8x8_stage_4_0_t101;
    FSM_dct_8x8_stage_4_0_t109[FSM_dct_8x8_stage_4_0_t104 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t108;
    FSM_dct_8x8_stage_4_0_t110 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_4_0_t111 = FSM_dct_8x8_stage_4_0_t110[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t112 = FSM_dct_8x8_stage_4_0_t111 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_4_0_t113 = FSM_dct_8x8_stage_4_0_t112[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t114 = FSM_dct_8x8_stage_4_0_t113[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t115 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_4_0_t116 = FSM_dct_8x8_stage_4_0_t115[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t117 = FSM_dct_8x8_stage_4_0_t116 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_4_0_t118 = FSM_dct_8x8_stage_4_0_t117[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t119 = FSM_dct_8x8_stage_4_0_t118[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t120 = i_data_in[FSM_dct_8x8_stage_4_0_t119 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t121 = FSM_dct_8x8_stage_4_0_t109;
    FSM_dct_8x8_stage_4_0_t121[FSM_dct_8x8_stage_4_0_t114 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t120;
    FSM_dct_8x8_stage_4_0_t122 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_4_0_t123 = FSM_dct_8x8_stage_4_0_t122[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t124 = FSM_dct_8x8_stage_4_0_t123 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_4_0_t125 = FSM_dct_8x8_stage_4_0_t124[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t126 = FSM_dct_8x8_stage_4_0_t125[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t127 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_4_0_t128 = FSM_dct_8x8_stage_4_0_t127[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t129 = FSM_dct_8x8_stage_4_0_t128 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_4_0_t130 = FSM_dct_8x8_stage_4_0_t129[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t131 = FSM_dct_8x8_stage_4_0_t130[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t132 = i_data_in[FSM_dct_8x8_stage_4_0_t131 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t133 = FSM_dct_8x8_stage_4_0_t132 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t134 = FSM_dct_8x8_stage_4_0_t133[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t135 = FSM_dct_8x8_stage_4_0_t121;
    FSM_dct_8x8_stage_4_0_t135[FSM_dct_8x8_stage_4_0_t126 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t134;
    FSM_dct_8x8_stage_4_0_t136 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_4_0_t137 = FSM_dct_8x8_stage_4_0_t136[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t138 = FSM_dct_8x8_stage_4_0_t137 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_4_0_t139 = FSM_dct_8x8_stage_4_0_t138[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t140 = FSM_dct_8x8_stage_4_0_t139[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t141 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_4_0_t142 = FSM_dct_8x8_stage_4_0_t141[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t143 = FSM_dct_8x8_stage_4_0_t142 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_4_0_t144 = FSM_dct_8x8_stage_4_0_t143[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t145 = FSM_dct_8x8_stage_4_0_t144[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t146 = i_data_in[FSM_dct_8x8_stage_4_0_t145 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t147 = FSM_dct_8x8_stage_4_0_t135;
    FSM_dct_8x8_stage_4_0_t147[FSM_dct_8x8_stage_4_0_t140 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t146;
    FSM_dct_8x8_stage_4_0_t148 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_4_0_t149 = FSM_dct_8x8_stage_4_0_t148[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t150 = FSM_dct_8x8_stage_4_0_t149 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_4_0_t151 = FSM_dct_8x8_stage_4_0_t150[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t152 = FSM_dct_8x8_stage_4_0_t151[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t153 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_4_0_t154 = FSM_dct_8x8_stage_4_0_t153[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t155 = FSM_dct_8x8_stage_4_0_t154 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_4_0_t156 = FSM_dct_8x8_stage_4_0_t155[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t157 = FSM_dct_8x8_stage_4_0_t156[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t158 = i_data_in[FSM_dct_8x8_stage_4_0_t157 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t159 = FSM_dct_8x8_stage_4_0_t158 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t160 = FSM_dct_8x8_stage_4_0_t159[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t161 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_4_0_t162 = FSM_dct_8x8_stage_4_0_t161[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t163 = FSM_dct_8x8_stage_4_0_t162 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_4_0_t164 = FSM_dct_8x8_stage_4_0_t163[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t165 = FSM_dct_8x8_stage_4_0_t164[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t166 = i_data_in[FSM_dct_8x8_stage_4_0_t165 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t167 = (FSM_dct_8x8_stage_4_0_t166 - FSM_dct_8x8_stage_4_0_t158) * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t168 = FSM_dct_8x8_stage_4_0_t167[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t169 = FSM_dct_8x8_stage_4_0_t147;
    FSM_dct_8x8_stage_4_0_t169[FSM_dct_8x8_stage_4_0_t152 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t160 - FSM_dct_8x8_stage_4_0_t168;
    FSM_dct_8x8_stage_4_0_t170 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_4_0_t171 = FSM_dct_8x8_stage_4_0_t170[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t172 = FSM_dct_8x8_stage_4_0_t171 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_4_0_t173 = FSM_dct_8x8_stage_4_0_t172[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t174 = FSM_dct_8x8_stage_4_0_t173[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t175 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_4_0_t176 = FSM_dct_8x8_stage_4_0_t175[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t177 = FSM_dct_8x8_stage_4_0_t176 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_4_0_t178 = FSM_dct_8x8_stage_4_0_t177[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t179 = FSM_dct_8x8_stage_4_0_t178[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t180 = i_data_in[FSM_dct_8x8_stage_4_0_t179 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t181 = FSM_dct_8x8_stage_4_0_t180 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t182 = FSM_dct_8x8_stage_4_0_t181[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t183 = FSM_dct_8x8_stage_4_0_t169;
    FSM_dct_8x8_stage_4_0_t183[FSM_dct_8x8_stage_4_0_t174 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t182;
    FSM_dct_8x8_stage_4_0_t184 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_4_0_t185 = FSM_dct_8x8_stage_4_0_t184[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t186 = FSM_dct_8x8_stage_4_0_t185 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_4_0_t187 = FSM_dct_8x8_stage_4_0_t186[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t188 = FSM_dct_8x8_stage_4_0_t187[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t189 = FSM_dct_8x8_stage_4_0_t166 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t190 = FSM_dct_8x8_stage_4_0_t189[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t191 = FSM_dct_8x8_stage_4_0_t183;
    FSM_dct_8x8_stage_4_0_t191[FSM_dct_8x8_stage_4_0_t188 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t190 - FSM_dct_8x8_stage_4_0_t168;
    FSM_dct_8x8_stage_4_0_t192 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_4_0_t193 = FSM_dct_8x8_stage_4_0_t192[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t194 = FSM_dct_8x8_stage_4_0_t193 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_4_0_t195 = FSM_dct_8x8_stage_4_0_t194[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t196 = FSM_dct_8x8_stage_4_0_t195[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t197 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_4_0_t198 = FSM_dct_8x8_stage_4_0_t197[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t199 = FSM_dct_8x8_stage_4_0_t198 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_4_0_t200 = FSM_dct_8x8_stage_4_0_t199[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t201 = FSM_dct_8x8_stage_4_0_t200[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t202 = i_data_in[FSM_dct_8x8_stage_4_0_t201 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t203 = FSM_dct_8x8_stage_4_0_t191;
    FSM_dct_8x8_stage_4_0_t203[FSM_dct_8x8_stage_4_0_t196 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t202;
    FSM_dct_8x8_stage_4_0_t204 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_4_0_t205 = FSM_dct_8x8_stage_4_0_t204[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t206 = FSM_dct_8x8_stage_4_0_t205[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t207 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_4_0_t208 = FSM_dct_8x8_stage_4_0_t207[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t209 = FSM_dct_8x8_stage_4_0_t208[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t210 = i_data_in[FSM_dct_8x8_stage_4_0_t209 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t211 = FSM_dct_8x8_stage_4_0_t203;
    FSM_dct_8x8_stage_4_0_t211[FSM_dct_8x8_stage_4_0_t206 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t210;
    FSM_dct_8x8_stage_4_0_t212 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_4_0_t213 = FSM_dct_8x8_stage_4_0_t212[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t214 = FSM_dct_8x8_stage_4_0_t213 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_4_0_t215 = FSM_dct_8x8_stage_4_0_t214[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t216 = FSM_dct_8x8_stage_4_0_t215[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t217 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_4_0_t218 = FSM_dct_8x8_stage_4_0_t217[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t219 = FSM_dct_8x8_stage_4_0_t218 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_4_0_t220 = FSM_dct_8x8_stage_4_0_t219[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t221 = FSM_dct_8x8_stage_4_0_t220[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t222 = i_data_in[FSM_dct_8x8_stage_4_0_t221 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t223 = FSM_dct_8x8_stage_4_0_t211;
    FSM_dct_8x8_stage_4_0_t223[FSM_dct_8x8_stage_4_0_t216 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t222;
    FSM_dct_8x8_stage_4_0_t224 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_4_0_t225 = FSM_dct_8x8_stage_4_0_t224[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t226 = FSM_dct_8x8_stage_4_0_t225 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_4_0_t227 = FSM_dct_8x8_stage_4_0_t226[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t228 = FSM_dct_8x8_stage_4_0_t227[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t229 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_4_0_t230 = FSM_dct_8x8_stage_4_0_t229[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t231 = FSM_dct_8x8_stage_4_0_t230 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_4_0_t232 = FSM_dct_8x8_stage_4_0_t231[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t233 = FSM_dct_8x8_stage_4_0_t232[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t234 = i_data_in[FSM_dct_8x8_stage_4_0_t233 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t235 = FSM_dct_8x8_stage_4_0_t234 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t236 = FSM_dct_8x8_stage_4_0_t235[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t237 = FSM_dct_8x8_stage_4_0_t223;
    FSM_dct_8x8_stage_4_0_t237[FSM_dct_8x8_stage_4_0_t228 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t236;
    FSM_dct_8x8_stage_4_0_t238 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_4_0_t239 = FSM_dct_8x8_stage_4_0_t238[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t240 = FSM_dct_8x8_stage_4_0_t239 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_4_0_t241 = FSM_dct_8x8_stage_4_0_t240[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t242 = FSM_dct_8x8_stage_4_0_t241[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t243 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_4_0_t244 = FSM_dct_8x8_stage_4_0_t243[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t245 = FSM_dct_8x8_stage_4_0_t244 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_4_0_t246 = FSM_dct_8x8_stage_4_0_t245[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t247 = FSM_dct_8x8_stage_4_0_t246[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t248 = i_data_in[FSM_dct_8x8_stage_4_0_t247 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t249 = FSM_dct_8x8_stage_4_0_t237;
    FSM_dct_8x8_stage_4_0_t249[FSM_dct_8x8_stage_4_0_t242 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t248;
    FSM_dct_8x8_stage_4_0_t250 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_4_0_t251 = FSM_dct_8x8_stage_4_0_t250[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t252 = FSM_dct_8x8_stage_4_0_t251 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_4_0_t253 = FSM_dct_8x8_stage_4_0_t252[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t254 = FSM_dct_8x8_stage_4_0_t253[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t255 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_4_0_t256 = FSM_dct_8x8_stage_4_0_t255[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t257 = FSM_dct_8x8_stage_4_0_t256 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_4_0_t258 = FSM_dct_8x8_stage_4_0_t257[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t259 = FSM_dct_8x8_stage_4_0_t258[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t260 = i_data_in[FSM_dct_8x8_stage_4_0_t259 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t261 = FSM_dct_8x8_stage_4_0_t260 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t262 = FSM_dct_8x8_stage_4_0_t261[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t263 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_4_0_t264 = FSM_dct_8x8_stage_4_0_t263[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t265 = FSM_dct_8x8_stage_4_0_t264 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_4_0_t266 = FSM_dct_8x8_stage_4_0_t265[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t267 = FSM_dct_8x8_stage_4_0_t266[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t268 = i_data_in[FSM_dct_8x8_stage_4_0_t267 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t269 = (FSM_dct_8x8_stage_4_0_t268 - FSM_dct_8x8_stage_4_0_t260) * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t270 = FSM_dct_8x8_stage_4_0_t269[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t271 = FSM_dct_8x8_stage_4_0_t249;
    FSM_dct_8x8_stage_4_0_t271[FSM_dct_8x8_stage_4_0_t254 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t262 - FSM_dct_8x8_stage_4_0_t270;
    FSM_dct_8x8_stage_4_0_t272 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_4_0_t273 = FSM_dct_8x8_stage_4_0_t272[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t274 = FSM_dct_8x8_stage_4_0_t273 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_4_0_t275 = FSM_dct_8x8_stage_4_0_t274[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t276 = FSM_dct_8x8_stage_4_0_t275[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t277 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_4_0_t278 = FSM_dct_8x8_stage_4_0_t277[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t279 = FSM_dct_8x8_stage_4_0_t278 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_4_0_t280 = FSM_dct_8x8_stage_4_0_t279[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t281 = FSM_dct_8x8_stage_4_0_t280[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t282 = i_data_in[FSM_dct_8x8_stage_4_0_t281 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t283 = FSM_dct_8x8_stage_4_0_t282 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t284 = FSM_dct_8x8_stage_4_0_t283[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t285 = FSM_dct_8x8_stage_4_0_t271;
    FSM_dct_8x8_stage_4_0_t285[FSM_dct_8x8_stage_4_0_t276 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t284;
    FSM_dct_8x8_stage_4_0_t286 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_4_0_t287 = FSM_dct_8x8_stage_4_0_t286[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t288 = FSM_dct_8x8_stage_4_0_t287 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_4_0_t289 = FSM_dct_8x8_stage_4_0_t288[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t290 = FSM_dct_8x8_stage_4_0_t289[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t291 = FSM_dct_8x8_stage_4_0_t268 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t292 = FSM_dct_8x8_stage_4_0_t291[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t293 = FSM_dct_8x8_stage_4_0_t285;
    FSM_dct_8x8_stage_4_0_t293[FSM_dct_8x8_stage_4_0_t290 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t292 - FSM_dct_8x8_stage_4_0_t270;
    FSM_dct_8x8_stage_4_0_t294 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_4_0_t295 = FSM_dct_8x8_stage_4_0_t294[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t296 = FSM_dct_8x8_stage_4_0_t295 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_4_0_t297 = FSM_dct_8x8_stage_4_0_t296[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t298 = FSM_dct_8x8_stage_4_0_t297[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t299 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_4_0_t300 = FSM_dct_8x8_stage_4_0_t299[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t301 = FSM_dct_8x8_stage_4_0_t300 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_4_0_t302 = FSM_dct_8x8_stage_4_0_t301[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t303 = FSM_dct_8x8_stage_4_0_t302[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t304 = i_data_in[FSM_dct_8x8_stage_4_0_t303 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t305 = FSM_dct_8x8_stage_4_0_t293;
    FSM_dct_8x8_stage_4_0_t305[FSM_dct_8x8_stage_4_0_t298 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t304;
    FSM_dct_8x8_stage_4_0_t306 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_4_0_t307 = FSM_dct_8x8_stage_4_0_t306[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t308 = FSM_dct_8x8_stage_4_0_t307[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t309 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_4_0_t310 = FSM_dct_8x8_stage_4_0_t309[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t311 = FSM_dct_8x8_stage_4_0_t310[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t312 = i_data_in[FSM_dct_8x8_stage_4_0_t311 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t313 = FSM_dct_8x8_stage_4_0_t305;
    FSM_dct_8x8_stage_4_0_t313[FSM_dct_8x8_stage_4_0_t308 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t312;
    FSM_dct_8x8_stage_4_0_t314 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_4_0_t315 = FSM_dct_8x8_stage_4_0_t314[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t316 = FSM_dct_8x8_stage_4_0_t315 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_4_0_t317 = FSM_dct_8x8_stage_4_0_t316[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t318 = FSM_dct_8x8_stage_4_0_t317[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t319 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_4_0_t320 = FSM_dct_8x8_stage_4_0_t319[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t321 = FSM_dct_8x8_stage_4_0_t320 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_4_0_t322 = FSM_dct_8x8_stage_4_0_t321[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t323 = FSM_dct_8x8_stage_4_0_t322[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t324 = i_data_in[FSM_dct_8x8_stage_4_0_t323 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t325 = FSM_dct_8x8_stage_4_0_t313;
    FSM_dct_8x8_stage_4_0_t325[FSM_dct_8x8_stage_4_0_t318 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t324;
    FSM_dct_8x8_stage_4_0_t326 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_4_0_t327 = FSM_dct_8x8_stage_4_0_t326[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t328 = FSM_dct_8x8_stage_4_0_t327 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_4_0_t329 = FSM_dct_8x8_stage_4_0_t328[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t330 = FSM_dct_8x8_stage_4_0_t329[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t331 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_4_0_t332 = FSM_dct_8x8_stage_4_0_t331[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t333 = FSM_dct_8x8_stage_4_0_t332 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_4_0_t334 = FSM_dct_8x8_stage_4_0_t333[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t335 = FSM_dct_8x8_stage_4_0_t334[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t336 = i_data_in[FSM_dct_8x8_stage_4_0_t335 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t337 = FSM_dct_8x8_stage_4_0_t336 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t338 = FSM_dct_8x8_stage_4_0_t337[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t339 = FSM_dct_8x8_stage_4_0_t325;
    FSM_dct_8x8_stage_4_0_t339[FSM_dct_8x8_stage_4_0_t330 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t338;
    FSM_dct_8x8_stage_4_0_t340 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_4_0_t341 = FSM_dct_8x8_stage_4_0_t340[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t342 = FSM_dct_8x8_stage_4_0_t341 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_4_0_t343 = FSM_dct_8x8_stage_4_0_t342[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t344 = FSM_dct_8x8_stage_4_0_t343[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t345 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_4_0_t346 = FSM_dct_8x8_stage_4_0_t345[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t347 = FSM_dct_8x8_stage_4_0_t346 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_4_0_t348 = FSM_dct_8x8_stage_4_0_t347[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t349 = FSM_dct_8x8_stage_4_0_t348[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t350 = i_data_in[FSM_dct_8x8_stage_4_0_t349 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t351 = FSM_dct_8x8_stage_4_0_t339;
    FSM_dct_8x8_stage_4_0_t351[FSM_dct_8x8_stage_4_0_t344 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t350;
    FSM_dct_8x8_stage_4_0_t352 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_4_0_t353 = FSM_dct_8x8_stage_4_0_t352[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t354 = FSM_dct_8x8_stage_4_0_t353 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_4_0_t355 = FSM_dct_8x8_stage_4_0_t354[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t356 = FSM_dct_8x8_stage_4_0_t355[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t357 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_4_0_t358 = FSM_dct_8x8_stage_4_0_t357[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t359 = FSM_dct_8x8_stage_4_0_t358 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_4_0_t360 = FSM_dct_8x8_stage_4_0_t359[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t361 = FSM_dct_8x8_stage_4_0_t360[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t362 = i_data_in[FSM_dct_8x8_stage_4_0_t361 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t363 = FSM_dct_8x8_stage_4_0_t362 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t364 = FSM_dct_8x8_stage_4_0_t363[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t365 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_4_0_t366 = FSM_dct_8x8_stage_4_0_t365[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t367 = FSM_dct_8x8_stage_4_0_t366 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_4_0_t368 = FSM_dct_8x8_stage_4_0_t367[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t369 = FSM_dct_8x8_stage_4_0_t368[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t370 = i_data_in[FSM_dct_8x8_stage_4_0_t369 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t371 = (FSM_dct_8x8_stage_4_0_t370 - FSM_dct_8x8_stage_4_0_t362) * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t372 = FSM_dct_8x8_stage_4_0_t371[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t373 = FSM_dct_8x8_stage_4_0_t351;
    FSM_dct_8x8_stage_4_0_t373[FSM_dct_8x8_stage_4_0_t356 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t364 - FSM_dct_8x8_stage_4_0_t372;
    FSM_dct_8x8_stage_4_0_t374 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_4_0_t375 = FSM_dct_8x8_stage_4_0_t374[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t376 = FSM_dct_8x8_stage_4_0_t375 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_4_0_t377 = FSM_dct_8x8_stage_4_0_t376[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t378 = FSM_dct_8x8_stage_4_0_t377[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t379 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_4_0_t380 = FSM_dct_8x8_stage_4_0_t379[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t381 = FSM_dct_8x8_stage_4_0_t380 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_4_0_t382 = FSM_dct_8x8_stage_4_0_t381[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t383 = FSM_dct_8x8_stage_4_0_t382[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t384 = i_data_in[FSM_dct_8x8_stage_4_0_t383 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t385 = FSM_dct_8x8_stage_4_0_t384 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t386 = FSM_dct_8x8_stage_4_0_t385[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t387 = FSM_dct_8x8_stage_4_0_t373;
    FSM_dct_8x8_stage_4_0_t387[FSM_dct_8x8_stage_4_0_t378 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t386;
    FSM_dct_8x8_stage_4_0_t388 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_4_0_t389 = FSM_dct_8x8_stage_4_0_t388[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t390 = FSM_dct_8x8_stage_4_0_t389 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_4_0_t391 = FSM_dct_8x8_stage_4_0_t390[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t392 = FSM_dct_8x8_stage_4_0_t391[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t393 = FSM_dct_8x8_stage_4_0_t370 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t394 = FSM_dct_8x8_stage_4_0_t393[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t395 = FSM_dct_8x8_stage_4_0_t387;
    FSM_dct_8x8_stage_4_0_t395[FSM_dct_8x8_stage_4_0_t392 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t394 - FSM_dct_8x8_stage_4_0_t372;
    FSM_dct_8x8_stage_4_0_t396 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_4_0_t397 = FSM_dct_8x8_stage_4_0_t396[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t398 = FSM_dct_8x8_stage_4_0_t397 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_4_0_t399 = FSM_dct_8x8_stage_4_0_t398[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t400 = FSM_dct_8x8_stage_4_0_t399[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t401 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_4_0_t402 = FSM_dct_8x8_stage_4_0_t401[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t403 = FSM_dct_8x8_stage_4_0_t402 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_4_0_t404 = FSM_dct_8x8_stage_4_0_t403[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t405 = FSM_dct_8x8_stage_4_0_t404[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t406 = i_data_in[FSM_dct_8x8_stage_4_0_t405 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t407 = FSM_dct_8x8_stage_4_0_t395;
    FSM_dct_8x8_stage_4_0_t407[FSM_dct_8x8_stage_4_0_t400 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t406;
    FSM_dct_8x8_stage_4_0_t408 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_4_0_t409 = FSM_dct_8x8_stage_4_0_t408[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t410 = FSM_dct_8x8_stage_4_0_t409[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t411 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_4_0_t412 = FSM_dct_8x8_stage_4_0_t411[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t413 = FSM_dct_8x8_stage_4_0_t412[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t414 = i_data_in[FSM_dct_8x8_stage_4_0_t413 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t415 = FSM_dct_8x8_stage_4_0_t407;
    FSM_dct_8x8_stage_4_0_t415[FSM_dct_8x8_stage_4_0_t410 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t414;
    FSM_dct_8x8_stage_4_0_t416 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_4_0_t417 = FSM_dct_8x8_stage_4_0_t416[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t418 = FSM_dct_8x8_stage_4_0_t417 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_4_0_t419 = FSM_dct_8x8_stage_4_0_t418[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t420 = FSM_dct_8x8_stage_4_0_t419[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t421 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_4_0_t422 = FSM_dct_8x8_stage_4_0_t421[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t423 = FSM_dct_8x8_stage_4_0_t422 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_4_0_t424 = FSM_dct_8x8_stage_4_0_t423[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t425 = FSM_dct_8x8_stage_4_0_t424[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t426 = i_data_in[FSM_dct_8x8_stage_4_0_t425 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t427 = FSM_dct_8x8_stage_4_0_t415;
    FSM_dct_8x8_stage_4_0_t427[FSM_dct_8x8_stage_4_0_t420 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t426;
    FSM_dct_8x8_stage_4_0_t428 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_4_0_t429 = FSM_dct_8x8_stage_4_0_t428[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t430 = FSM_dct_8x8_stage_4_0_t429 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_4_0_t431 = FSM_dct_8x8_stage_4_0_t430[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t432 = FSM_dct_8x8_stage_4_0_t431[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t433 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_4_0_t434 = FSM_dct_8x8_stage_4_0_t433[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t435 = FSM_dct_8x8_stage_4_0_t434 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_4_0_t436 = FSM_dct_8x8_stage_4_0_t435[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t437 = FSM_dct_8x8_stage_4_0_t436[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t438 = i_data_in[FSM_dct_8x8_stage_4_0_t437 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t439 = FSM_dct_8x8_stage_4_0_t438 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t440 = FSM_dct_8x8_stage_4_0_t439[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t441 = FSM_dct_8x8_stage_4_0_t427;
    FSM_dct_8x8_stage_4_0_t441[FSM_dct_8x8_stage_4_0_t432 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t440;
    FSM_dct_8x8_stage_4_0_t442 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_4_0_t443 = FSM_dct_8x8_stage_4_0_t442[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t444 = FSM_dct_8x8_stage_4_0_t443 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_4_0_t445 = FSM_dct_8x8_stage_4_0_t444[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t446 = FSM_dct_8x8_stage_4_0_t445[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t447 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_4_0_t448 = FSM_dct_8x8_stage_4_0_t447[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t449 = FSM_dct_8x8_stage_4_0_t448 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_4_0_t450 = FSM_dct_8x8_stage_4_0_t449[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t451 = FSM_dct_8x8_stage_4_0_t450[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t452 = i_data_in[FSM_dct_8x8_stage_4_0_t451 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t453 = FSM_dct_8x8_stage_4_0_t441;
    FSM_dct_8x8_stage_4_0_t453[FSM_dct_8x8_stage_4_0_t446 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t452;
    FSM_dct_8x8_stage_4_0_t454 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_4_0_t455 = FSM_dct_8x8_stage_4_0_t454[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t456 = FSM_dct_8x8_stage_4_0_t455 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_4_0_t457 = FSM_dct_8x8_stage_4_0_t456[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t458 = FSM_dct_8x8_stage_4_0_t457[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t459 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_4_0_t460 = FSM_dct_8x8_stage_4_0_t459[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t461 = FSM_dct_8x8_stage_4_0_t460 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_4_0_t462 = FSM_dct_8x8_stage_4_0_t461[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t463 = FSM_dct_8x8_stage_4_0_t462[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t464 = i_data_in[FSM_dct_8x8_stage_4_0_t463 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t465 = FSM_dct_8x8_stage_4_0_t464 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t466 = FSM_dct_8x8_stage_4_0_t465[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t467 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_4_0_t468 = FSM_dct_8x8_stage_4_0_t467[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t469 = FSM_dct_8x8_stage_4_0_t468 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_4_0_t470 = FSM_dct_8x8_stage_4_0_t469[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t471 = FSM_dct_8x8_stage_4_0_t470[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t472 = i_data_in[FSM_dct_8x8_stage_4_0_t471 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t473 = (FSM_dct_8x8_stage_4_0_t472 - FSM_dct_8x8_stage_4_0_t464) * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t474 = FSM_dct_8x8_stage_4_0_t473[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t475 = FSM_dct_8x8_stage_4_0_t453;
    FSM_dct_8x8_stage_4_0_t475[FSM_dct_8x8_stage_4_0_t458 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t466 - FSM_dct_8x8_stage_4_0_t474;
    FSM_dct_8x8_stage_4_0_t476 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_4_0_t477 = FSM_dct_8x8_stage_4_0_t476[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t478 = FSM_dct_8x8_stage_4_0_t477 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_4_0_t479 = FSM_dct_8x8_stage_4_0_t478[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t480 = FSM_dct_8x8_stage_4_0_t479[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t481 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_4_0_t482 = FSM_dct_8x8_stage_4_0_t481[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t483 = FSM_dct_8x8_stage_4_0_t482 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_4_0_t484 = FSM_dct_8x8_stage_4_0_t483[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t485 = FSM_dct_8x8_stage_4_0_t484[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t486 = i_data_in[FSM_dct_8x8_stage_4_0_t485 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t487 = FSM_dct_8x8_stage_4_0_t486 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t488 = FSM_dct_8x8_stage_4_0_t487[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t489 = FSM_dct_8x8_stage_4_0_t475;
    FSM_dct_8x8_stage_4_0_t489[FSM_dct_8x8_stage_4_0_t480 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t488;
    FSM_dct_8x8_stage_4_0_t490 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_4_0_t491 = FSM_dct_8x8_stage_4_0_t490[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t492 = FSM_dct_8x8_stage_4_0_t491 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_4_0_t493 = FSM_dct_8x8_stage_4_0_t492[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t494 = FSM_dct_8x8_stage_4_0_t493[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t495 = FSM_dct_8x8_stage_4_0_t472 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t496 = FSM_dct_8x8_stage_4_0_t495[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t497 = FSM_dct_8x8_stage_4_0_t489;
    FSM_dct_8x8_stage_4_0_t497[FSM_dct_8x8_stage_4_0_t494 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t496 - FSM_dct_8x8_stage_4_0_t474;
    FSM_dct_8x8_stage_4_0_t498 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_4_0_t499 = FSM_dct_8x8_stage_4_0_t498[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t500 = FSM_dct_8x8_stage_4_0_t499 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_4_0_t501 = FSM_dct_8x8_stage_4_0_t500[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t502 = FSM_dct_8x8_stage_4_0_t501[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t503 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_4_0_t504 = FSM_dct_8x8_stage_4_0_t503[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t505 = FSM_dct_8x8_stage_4_0_t504 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_4_0_t506 = FSM_dct_8x8_stage_4_0_t505[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t507 = FSM_dct_8x8_stage_4_0_t506[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t508 = i_data_in[FSM_dct_8x8_stage_4_0_t507 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t509 = FSM_dct_8x8_stage_4_0_t497;
    FSM_dct_8x8_stage_4_0_t509[FSM_dct_8x8_stage_4_0_t502 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t508;
    FSM_dct_8x8_stage_4_0_t510 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_4_0_t511 = FSM_dct_8x8_stage_4_0_t510[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t512 = FSM_dct_8x8_stage_4_0_t511[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t513 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_4_0_t514 = FSM_dct_8x8_stage_4_0_t513[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t515 = FSM_dct_8x8_stage_4_0_t514[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t516 = i_data_in[FSM_dct_8x8_stage_4_0_t515 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t517 = FSM_dct_8x8_stage_4_0_t509;
    FSM_dct_8x8_stage_4_0_t517[FSM_dct_8x8_stage_4_0_t512 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t516;
    FSM_dct_8x8_stage_4_0_t518 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_4_0_t519 = FSM_dct_8x8_stage_4_0_t518[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t520 = FSM_dct_8x8_stage_4_0_t519 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_4_0_t521 = FSM_dct_8x8_stage_4_0_t520[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t522 = FSM_dct_8x8_stage_4_0_t521[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t523 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_4_0_t524 = FSM_dct_8x8_stage_4_0_t523[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t525 = FSM_dct_8x8_stage_4_0_t524 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_4_0_t526 = FSM_dct_8x8_stage_4_0_t525[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t527 = FSM_dct_8x8_stage_4_0_t526[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t528 = i_data_in[FSM_dct_8x8_stage_4_0_t527 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t529 = FSM_dct_8x8_stage_4_0_t517;
    FSM_dct_8x8_stage_4_0_t529[FSM_dct_8x8_stage_4_0_t522 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t528;
    FSM_dct_8x8_stage_4_0_t530 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_4_0_t531 = FSM_dct_8x8_stage_4_0_t530[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t532 = FSM_dct_8x8_stage_4_0_t531 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_4_0_t533 = FSM_dct_8x8_stage_4_0_t532[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t534 = FSM_dct_8x8_stage_4_0_t533[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t535 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_4_0_t536 = FSM_dct_8x8_stage_4_0_t535[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t537 = FSM_dct_8x8_stage_4_0_t536 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_4_0_t538 = FSM_dct_8x8_stage_4_0_t537[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t539 = FSM_dct_8x8_stage_4_0_t538[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t540 = i_data_in[FSM_dct_8x8_stage_4_0_t539 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t541 = FSM_dct_8x8_stage_4_0_t540 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t542 = FSM_dct_8x8_stage_4_0_t541[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t543 = FSM_dct_8x8_stage_4_0_t529;
    FSM_dct_8x8_stage_4_0_t543[FSM_dct_8x8_stage_4_0_t534 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t542;
    FSM_dct_8x8_stage_4_0_t544 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_4_0_t545 = FSM_dct_8x8_stage_4_0_t544[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t546 = FSM_dct_8x8_stage_4_0_t545 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_4_0_t547 = FSM_dct_8x8_stage_4_0_t546[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t548 = FSM_dct_8x8_stage_4_0_t547[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t549 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_4_0_t550 = FSM_dct_8x8_stage_4_0_t549[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t551 = FSM_dct_8x8_stage_4_0_t550 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_4_0_t552 = FSM_dct_8x8_stage_4_0_t551[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t553 = FSM_dct_8x8_stage_4_0_t552[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t554 = i_data_in[FSM_dct_8x8_stage_4_0_t553 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t555 = FSM_dct_8x8_stage_4_0_t543;
    FSM_dct_8x8_stage_4_0_t555[FSM_dct_8x8_stage_4_0_t548 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t554;
    FSM_dct_8x8_stage_4_0_t556 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_4_0_t557 = FSM_dct_8x8_stage_4_0_t556[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t558 = FSM_dct_8x8_stage_4_0_t557 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_4_0_t559 = FSM_dct_8x8_stage_4_0_t558[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t560 = FSM_dct_8x8_stage_4_0_t559[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t561 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_4_0_t562 = FSM_dct_8x8_stage_4_0_t561[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t563 = FSM_dct_8x8_stage_4_0_t562 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_4_0_t564 = FSM_dct_8x8_stage_4_0_t563[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t565 = FSM_dct_8x8_stage_4_0_t564[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t566 = i_data_in[FSM_dct_8x8_stage_4_0_t565 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t567 = FSM_dct_8x8_stage_4_0_t566 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t568 = FSM_dct_8x8_stage_4_0_t567[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t569 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_4_0_t570 = FSM_dct_8x8_stage_4_0_t569[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t571 = FSM_dct_8x8_stage_4_0_t570 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_4_0_t572 = FSM_dct_8x8_stage_4_0_t571[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t573 = FSM_dct_8x8_stage_4_0_t572[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t574 = i_data_in[FSM_dct_8x8_stage_4_0_t573 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t575 = (FSM_dct_8x8_stage_4_0_t574 - FSM_dct_8x8_stage_4_0_t566) * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t576 = FSM_dct_8x8_stage_4_0_t575[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t577 = FSM_dct_8x8_stage_4_0_t555;
    FSM_dct_8x8_stage_4_0_t577[FSM_dct_8x8_stage_4_0_t560 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t568 - FSM_dct_8x8_stage_4_0_t576;
    FSM_dct_8x8_stage_4_0_t578 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_4_0_t579 = FSM_dct_8x8_stage_4_0_t578[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t580 = FSM_dct_8x8_stage_4_0_t579 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_4_0_t581 = FSM_dct_8x8_stage_4_0_t580[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t582 = FSM_dct_8x8_stage_4_0_t581[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t583 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_4_0_t584 = FSM_dct_8x8_stage_4_0_t583[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t585 = FSM_dct_8x8_stage_4_0_t584 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_4_0_t586 = FSM_dct_8x8_stage_4_0_t585[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t587 = FSM_dct_8x8_stage_4_0_t586[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t588 = i_data_in[FSM_dct_8x8_stage_4_0_t587 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t589 = FSM_dct_8x8_stage_4_0_t588 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t590 = FSM_dct_8x8_stage_4_0_t589[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t591 = FSM_dct_8x8_stage_4_0_t577;
    FSM_dct_8x8_stage_4_0_t591[FSM_dct_8x8_stage_4_0_t582 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t590;
    FSM_dct_8x8_stage_4_0_t592 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_4_0_t593 = FSM_dct_8x8_stage_4_0_t592[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t594 = FSM_dct_8x8_stage_4_0_t593 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_4_0_t595 = FSM_dct_8x8_stage_4_0_t594[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t596 = FSM_dct_8x8_stage_4_0_t595[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t597 = FSM_dct_8x8_stage_4_0_t574 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t598 = FSM_dct_8x8_stage_4_0_t597[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t599 = FSM_dct_8x8_stage_4_0_t591;
    FSM_dct_8x8_stage_4_0_t599[FSM_dct_8x8_stage_4_0_t596 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t598 - FSM_dct_8x8_stage_4_0_t576;
    FSM_dct_8x8_stage_4_0_t600 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_4_0_t601 = FSM_dct_8x8_stage_4_0_t600[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t602 = FSM_dct_8x8_stage_4_0_t601 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_4_0_t603 = FSM_dct_8x8_stage_4_0_t602[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t604 = FSM_dct_8x8_stage_4_0_t603[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t605 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_4_0_t606 = FSM_dct_8x8_stage_4_0_t605[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t607 = FSM_dct_8x8_stage_4_0_t606 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_4_0_t608 = FSM_dct_8x8_stage_4_0_t607[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t609 = FSM_dct_8x8_stage_4_0_t608[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t610 = i_data_in[FSM_dct_8x8_stage_4_0_t609 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t611 = FSM_dct_8x8_stage_4_0_t599;
    FSM_dct_8x8_stage_4_0_t611[FSM_dct_8x8_stage_4_0_t604 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t610;
    FSM_dct_8x8_stage_4_0_t612 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_4_0_t613 = FSM_dct_8x8_stage_4_0_t612[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t614 = FSM_dct_8x8_stage_4_0_t613[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t615 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_4_0_t616 = FSM_dct_8x8_stage_4_0_t615[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t617 = FSM_dct_8x8_stage_4_0_t616[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t618 = i_data_in[FSM_dct_8x8_stage_4_0_t617 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t619 = FSM_dct_8x8_stage_4_0_t611;
    FSM_dct_8x8_stage_4_0_t619[FSM_dct_8x8_stage_4_0_t614 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t618;
    FSM_dct_8x8_stage_4_0_t620 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_4_0_t621 = FSM_dct_8x8_stage_4_0_t620[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t622 = FSM_dct_8x8_stage_4_0_t621 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_4_0_t623 = FSM_dct_8x8_stage_4_0_t622[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t624 = FSM_dct_8x8_stage_4_0_t623[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t625 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_4_0_t626 = FSM_dct_8x8_stage_4_0_t625[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t627 = FSM_dct_8x8_stage_4_0_t626 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_4_0_t628 = FSM_dct_8x8_stage_4_0_t627[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t629 = FSM_dct_8x8_stage_4_0_t628[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t630 = i_data_in[FSM_dct_8x8_stage_4_0_t629 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t631 = FSM_dct_8x8_stage_4_0_t619;
    FSM_dct_8x8_stage_4_0_t631[FSM_dct_8x8_stage_4_0_t624 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t630;
    FSM_dct_8x8_stage_4_0_t632 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_4_0_t633 = FSM_dct_8x8_stage_4_0_t632[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t634 = FSM_dct_8x8_stage_4_0_t633 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_4_0_t635 = FSM_dct_8x8_stage_4_0_t634[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t636 = FSM_dct_8x8_stage_4_0_t635[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t637 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_4_0_t638 = FSM_dct_8x8_stage_4_0_t637[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t639 = FSM_dct_8x8_stage_4_0_t638 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_4_0_t640 = FSM_dct_8x8_stage_4_0_t639[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t641 = FSM_dct_8x8_stage_4_0_t640[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t642 = i_data_in[FSM_dct_8x8_stage_4_0_t641 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t643 = FSM_dct_8x8_stage_4_0_t642 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t644 = FSM_dct_8x8_stage_4_0_t643[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t645 = FSM_dct_8x8_stage_4_0_t631;
    FSM_dct_8x8_stage_4_0_t645[FSM_dct_8x8_stage_4_0_t636 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t644;
    FSM_dct_8x8_stage_4_0_t646 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_4_0_t647 = FSM_dct_8x8_stage_4_0_t646[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t648 = FSM_dct_8x8_stage_4_0_t647 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_4_0_t649 = FSM_dct_8x8_stage_4_0_t648[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t650 = FSM_dct_8x8_stage_4_0_t649[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t651 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_4_0_t652 = FSM_dct_8x8_stage_4_0_t651[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t653 = FSM_dct_8x8_stage_4_0_t652 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_4_0_t654 = FSM_dct_8x8_stage_4_0_t653[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t655 = FSM_dct_8x8_stage_4_0_t654[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t656 = i_data_in[FSM_dct_8x8_stage_4_0_t655 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t657 = FSM_dct_8x8_stage_4_0_t645;
    FSM_dct_8x8_stage_4_0_t657[FSM_dct_8x8_stage_4_0_t650 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t656;
    FSM_dct_8x8_stage_4_0_t658 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_4_0_t659 = FSM_dct_8x8_stage_4_0_t658[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t660 = FSM_dct_8x8_stage_4_0_t659 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_4_0_t661 = FSM_dct_8x8_stage_4_0_t660[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t662 = FSM_dct_8x8_stage_4_0_t661[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t663 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_4_0_t664 = FSM_dct_8x8_stage_4_0_t663[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t665 = FSM_dct_8x8_stage_4_0_t664 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_4_0_t666 = FSM_dct_8x8_stage_4_0_t665[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t667 = FSM_dct_8x8_stage_4_0_t666[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t668 = i_data_in[FSM_dct_8x8_stage_4_0_t667 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t669 = FSM_dct_8x8_stage_4_0_t668 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t670 = FSM_dct_8x8_stage_4_0_t669[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t671 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_4_0_t672 = FSM_dct_8x8_stage_4_0_t671[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t673 = FSM_dct_8x8_stage_4_0_t672 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_4_0_t674 = FSM_dct_8x8_stage_4_0_t673[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t675 = FSM_dct_8x8_stage_4_0_t674[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t676 = i_data_in[FSM_dct_8x8_stage_4_0_t675 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t677 = (FSM_dct_8x8_stage_4_0_t676 - FSM_dct_8x8_stage_4_0_t668) * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t678 = FSM_dct_8x8_stage_4_0_t677[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t679 = FSM_dct_8x8_stage_4_0_t657;
    FSM_dct_8x8_stage_4_0_t679[FSM_dct_8x8_stage_4_0_t662 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t670 - FSM_dct_8x8_stage_4_0_t678;
    FSM_dct_8x8_stage_4_0_t680 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_4_0_t681 = FSM_dct_8x8_stage_4_0_t680[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t682 = FSM_dct_8x8_stage_4_0_t681 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_4_0_t683 = FSM_dct_8x8_stage_4_0_t682[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t684 = FSM_dct_8x8_stage_4_0_t683[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t685 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_4_0_t686 = FSM_dct_8x8_stage_4_0_t685[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t687 = FSM_dct_8x8_stage_4_0_t686 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_4_0_t688 = FSM_dct_8x8_stage_4_0_t687[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t689 = FSM_dct_8x8_stage_4_0_t688[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t690 = i_data_in[FSM_dct_8x8_stage_4_0_t689 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t691 = FSM_dct_8x8_stage_4_0_t690 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t692 = FSM_dct_8x8_stage_4_0_t691[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t693 = FSM_dct_8x8_stage_4_0_t679;
    FSM_dct_8x8_stage_4_0_t693[FSM_dct_8x8_stage_4_0_t684 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t692;
    FSM_dct_8x8_stage_4_0_t694 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_4_0_t695 = FSM_dct_8x8_stage_4_0_t694[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t696 = FSM_dct_8x8_stage_4_0_t695 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_4_0_t697 = FSM_dct_8x8_stage_4_0_t696[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t698 = FSM_dct_8x8_stage_4_0_t697[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t699 = FSM_dct_8x8_stage_4_0_t676 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t700 = FSM_dct_8x8_stage_4_0_t699[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t701 = FSM_dct_8x8_stage_4_0_t693;
    FSM_dct_8x8_stage_4_0_t701[FSM_dct_8x8_stage_4_0_t698 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t700 - FSM_dct_8x8_stage_4_0_t678;
    FSM_dct_8x8_stage_4_0_t702 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_4_0_t703 = FSM_dct_8x8_stage_4_0_t702[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t704 = FSM_dct_8x8_stage_4_0_t703 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_4_0_t705 = FSM_dct_8x8_stage_4_0_t704[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t706 = FSM_dct_8x8_stage_4_0_t705[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t707 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_4_0_t708 = FSM_dct_8x8_stage_4_0_t707[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t709 = FSM_dct_8x8_stage_4_0_t708 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_4_0_t710 = FSM_dct_8x8_stage_4_0_t709[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t711 = FSM_dct_8x8_stage_4_0_t710[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t712 = i_data_in[FSM_dct_8x8_stage_4_0_t711 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t713 = FSM_dct_8x8_stage_4_0_t701;
    FSM_dct_8x8_stage_4_0_t713[FSM_dct_8x8_stage_4_0_t706 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t712;
    FSM_dct_8x8_stage_4_0_t714 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_4_0_t715 = FSM_dct_8x8_stage_4_0_t714[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t716 = FSM_dct_8x8_stage_4_0_t715[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t717 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_4_0_t718 = FSM_dct_8x8_stage_4_0_t717[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t719 = FSM_dct_8x8_stage_4_0_t718[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t720 = i_data_in[FSM_dct_8x8_stage_4_0_t719 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t721 = FSM_dct_8x8_stage_4_0_t713;
    FSM_dct_8x8_stage_4_0_t721[FSM_dct_8x8_stage_4_0_t716 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t720;
    FSM_dct_8x8_stage_4_0_t722 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_4_0_t723 = FSM_dct_8x8_stage_4_0_t722[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t724 = FSM_dct_8x8_stage_4_0_t723 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_4_0_t725 = FSM_dct_8x8_stage_4_0_t724[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t726 = FSM_dct_8x8_stage_4_0_t725[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t727 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_4_0_t728 = FSM_dct_8x8_stage_4_0_t727[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t729 = FSM_dct_8x8_stage_4_0_t728 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_4_0_t730 = FSM_dct_8x8_stage_4_0_t729[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t731 = FSM_dct_8x8_stage_4_0_t730[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t732 = i_data_in[FSM_dct_8x8_stage_4_0_t731 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t733 = FSM_dct_8x8_stage_4_0_t721;
    FSM_dct_8x8_stage_4_0_t733[FSM_dct_8x8_stage_4_0_t726 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t732;
    FSM_dct_8x8_stage_4_0_t734 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_4_0_t735 = FSM_dct_8x8_stage_4_0_t734[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t736 = FSM_dct_8x8_stage_4_0_t735 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_4_0_t737 = FSM_dct_8x8_stage_4_0_t736[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t738 = FSM_dct_8x8_stage_4_0_t737[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t739 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_4_0_t740 = FSM_dct_8x8_stage_4_0_t739[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t741 = FSM_dct_8x8_stage_4_0_t740 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_4_0_t742 = FSM_dct_8x8_stage_4_0_t741[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t743 = FSM_dct_8x8_stage_4_0_t742[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t744 = i_data_in[FSM_dct_8x8_stage_4_0_t743 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t745 = FSM_dct_8x8_stage_4_0_t744 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t746 = FSM_dct_8x8_stage_4_0_t745[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t747 = FSM_dct_8x8_stage_4_0_t733;
    FSM_dct_8x8_stage_4_0_t747[FSM_dct_8x8_stage_4_0_t738 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t746;
    FSM_dct_8x8_stage_4_0_t748 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_4_0_t749 = FSM_dct_8x8_stage_4_0_t748[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t750 = FSM_dct_8x8_stage_4_0_t749 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_4_0_t751 = FSM_dct_8x8_stage_4_0_t750[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t752 = FSM_dct_8x8_stage_4_0_t751[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t753 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_4_0_t754 = FSM_dct_8x8_stage_4_0_t753[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t755 = FSM_dct_8x8_stage_4_0_t754 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_4_0_t756 = FSM_dct_8x8_stage_4_0_t755[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t757 = FSM_dct_8x8_stage_4_0_t756[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t758 = i_data_in[FSM_dct_8x8_stage_4_0_t757 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t759 = FSM_dct_8x8_stage_4_0_t747;
    FSM_dct_8x8_stage_4_0_t759[FSM_dct_8x8_stage_4_0_t752 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t758;
    FSM_dct_8x8_stage_4_0_t760 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_4_0_t761 = FSM_dct_8x8_stage_4_0_t760[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t762 = FSM_dct_8x8_stage_4_0_t761 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_4_0_t763 = FSM_dct_8x8_stage_4_0_t762[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t764 = FSM_dct_8x8_stage_4_0_t763[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t765 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_4_0_t766 = FSM_dct_8x8_stage_4_0_t765[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t767 = FSM_dct_8x8_stage_4_0_t766 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_4_0_t768 = FSM_dct_8x8_stage_4_0_t767[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t769 = FSM_dct_8x8_stage_4_0_t768[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t770 = i_data_in[FSM_dct_8x8_stage_4_0_t769 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t771 = FSM_dct_8x8_stage_4_0_t770 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t772 = FSM_dct_8x8_stage_4_0_t771[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t773 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_4_0_t774 = FSM_dct_8x8_stage_4_0_t773[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t775 = FSM_dct_8x8_stage_4_0_t774 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_4_0_t776 = FSM_dct_8x8_stage_4_0_t775[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t777 = FSM_dct_8x8_stage_4_0_t776[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t778 = i_data_in[FSM_dct_8x8_stage_4_0_t777 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t779 = (FSM_dct_8x8_stage_4_0_t778 - FSM_dct_8x8_stage_4_0_t770) * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t780 = FSM_dct_8x8_stage_4_0_t779[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t781 = FSM_dct_8x8_stage_4_0_t759;
    FSM_dct_8x8_stage_4_0_t781[FSM_dct_8x8_stage_4_0_t764 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t772 - FSM_dct_8x8_stage_4_0_t780;
    FSM_dct_8x8_stage_4_0_t782 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_4_0_t783 = FSM_dct_8x8_stage_4_0_t782[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t784 = FSM_dct_8x8_stage_4_0_t783 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_4_0_t785 = FSM_dct_8x8_stage_4_0_t784[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t786 = FSM_dct_8x8_stage_4_0_t785[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t787 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_4_0_t788 = FSM_dct_8x8_stage_4_0_t787[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t789 = FSM_dct_8x8_stage_4_0_t788 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_4_0_t790 = FSM_dct_8x8_stage_4_0_t789[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t791 = FSM_dct_8x8_stage_4_0_t790[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t792 = i_data_in[FSM_dct_8x8_stage_4_0_t791 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t793 = FSM_dct_8x8_stage_4_0_t792 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t794 = FSM_dct_8x8_stage_4_0_t793[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t795 = FSM_dct_8x8_stage_4_0_t781;
    FSM_dct_8x8_stage_4_0_t795[FSM_dct_8x8_stage_4_0_t786 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t794;
    FSM_dct_8x8_stage_4_0_t796 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_4_0_t797 = FSM_dct_8x8_stage_4_0_t796[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t798 = FSM_dct_8x8_stage_4_0_t797 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_4_0_t799 = FSM_dct_8x8_stage_4_0_t798[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t800 = FSM_dct_8x8_stage_4_0_t799[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t801 = FSM_dct_8x8_stage_4_0_t778 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t802 = FSM_dct_8x8_stage_4_0_t801[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t803 = FSM_dct_8x8_stage_4_0_t795;
    FSM_dct_8x8_stage_4_0_t803[FSM_dct_8x8_stage_4_0_t800 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t802 - FSM_dct_8x8_stage_4_0_t780;
    FSM_dct_8x8_stage_4_0_t804 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_4_0_t805 = FSM_dct_8x8_stage_4_0_t804[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t806 = FSM_dct_8x8_stage_4_0_t805 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_4_0_t807 = FSM_dct_8x8_stage_4_0_t806[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t808 = FSM_dct_8x8_stage_4_0_t807[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t809 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_4_0_t810 = FSM_dct_8x8_stage_4_0_t809[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t811 = FSM_dct_8x8_stage_4_0_t810 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_4_0_t812 = FSM_dct_8x8_stage_4_0_t811[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t813 = FSM_dct_8x8_stage_4_0_t812[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t814 = i_data_in[FSM_dct_8x8_stage_4_0_t813 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t815 = FSM_dct_8x8_stage_4_0_t803;
    FSM_dct_8x8_stage_4_0_t815[FSM_dct_8x8_stage_4_0_t808 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t814;
end

always @* begin
    FSM_dct_8x8_stage_4_0_t0 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_4_0_t1 = FSM_dct_8x8_stage_4_0_t0[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t2 = FSM_dct_8x8_stage_4_0_t1[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t3 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_4_0_t4 = FSM_dct_8x8_stage_4_0_t3[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t5 = FSM_dct_8x8_stage_4_0_t4[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t6 = i_data_in[FSM_dct_8x8_stage_4_0_t5 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t7 = 2048'b0;
    FSM_dct_8x8_stage_4_0_t7[FSM_dct_8x8_stage_4_0_t2 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t6;
    FSM_dct_8x8_stage_4_0_t8 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_4_0_t9 = FSM_dct_8x8_stage_4_0_t8[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t10 = FSM_dct_8x8_stage_4_0_t9 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_4_0_t11 = FSM_dct_8x8_stage_4_0_t10[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t12 = FSM_dct_8x8_stage_4_0_t11[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t13 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_4_0_t14 = FSM_dct_8x8_stage_4_0_t13[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t15 = FSM_dct_8x8_stage_4_0_t14 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_4_0_t16 = FSM_dct_8x8_stage_4_0_t15[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t17 = FSM_dct_8x8_stage_4_0_t16[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t18 = i_data_in[FSM_dct_8x8_stage_4_0_t17 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t19 = FSM_dct_8x8_stage_4_0_t7;
    FSM_dct_8x8_stage_4_0_t19[FSM_dct_8x8_stage_4_0_t12 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t18;
    FSM_dct_8x8_stage_4_0_t20 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_4_0_t21 = FSM_dct_8x8_stage_4_0_t20[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t22 = FSM_dct_8x8_stage_4_0_t21 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_4_0_t23 = FSM_dct_8x8_stage_4_0_t22[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t24 = FSM_dct_8x8_stage_4_0_t23[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t25 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_4_0_t26 = FSM_dct_8x8_stage_4_0_t25[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t27 = FSM_dct_8x8_stage_4_0_t26 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_4_0_t28 = FSM_dct_8x8_stage_4_0_t27[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t29 = FSM_dct_8x8_stage_4_0_t28[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t30 = i_data_in[FSM_dct_8x8_stage_4_0_t29 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t31 = FSM_dct_8x8_stage_4_0_t30 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t32 = FSM_dct_8x8_stage_4_0_t31[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t33 = FSM_dct_8x8_stage_4_0_t19;
    FSM_dct_8x8_stage_4_0_t33[FSM_dct_8x8_stage_4_0_t24 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t32;
    FSM_dct_8x8_stage_4_0_t34 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_4_0_t35 = FSM_dct_8x8_stage_4_0_t34[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t36 = FSM_dct_8x8_stage_4_0_t35 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_4_0_t37 = FSM_dct_8x8_stage_4_0_t36[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t38 = FSM_dct_8x8_stage_4_0_t37[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t39 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_4_0_t40 = FSM_dct_8x8_stage_4_0_t39[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t41 = FSM_dct_8x8_stage_4_0_t40 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_4_0_t42 = FSM_dct_8x8_stage_4_0_t41[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t43 = FSM_dct_8x8_stage_4_0_t42[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t44 = i_data_in[FSM_dct_8x8_stage_4_0_t43 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t45 = FSM_dct_8x8_stage_4_0_t33;
    FSM_dct_8x8_stage_4_0_t45[FSM_dct_8x8_stage_4_0_t38 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t44;
    FSM_dct_8x8_stage_4_0_t46 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_4_0_t47 = FSM_dct_8x8_stage_4_0_t46[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t48 = FSM_dct_8x8_stage_4_0_t47 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_4_0_t49 = FSM_dct_8x8_stage_4_0_t48[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t50 = FSM_dct_8x8_stage_4_0_t49[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t51 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_4_0_t52 = FSM_dct_8x8_stage_4_0_t51[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t53 = FSM_dct_8x8_stage_4_0_t52 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_4_0_t54 = FSM_dct_8x8_stage_4_0_t53[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t55 = FSM_dct_8x8_stage_4_0_t54[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t56 = i_data_in[FSM_dct_8x8_stage_4_0_t55 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t57 = FSM_dct_8x8_stage_4_0_t56 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t58 = FSM_dct_8x8_stage_4_0_t57[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t59 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_4_0_t60 = FSM_dct_8x8_stage_4_0_t59[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t61 = FSM_dct_8x8_stage_4_0_t60 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_4_0_t62 = FSM_dct_8x8_stage_4_0_t61[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t63 = FSM_dct_8x8_stage_4_0_t62[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t64 = i_data_in[FSM_dct_8x8_stage_4_0_t63 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t65 = (FSM_dct_8x8_stage_4_0_t64 - FSM_dct_8x8_stage_4_0_t56) * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t66 = FSM_dct_8x8_stage_4_0_t65[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t67 = FSM_dct_8x8_stage_4_0_t45;
    FSM_dct_8x8_stage_4_0_t67[FSM_dct_8x8_stage_4_0_t50 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t58 - FSM_dct_8x8_stage_4_0_t66;
    FSM_dct_8x8_stage_4_0_t68 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_4_0_t69 = FSM_dct_8x8_stage_4_0_t68[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t70 = FSM_dct_8x8_stage_4_0_t69 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_4_0_t71 = FSM_dct_8x8_stage_4_0_t70[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t72 = FSM_dct_8x8_stage_4_0_t71[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t73 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_4_0_t74 = FSM_dct_8x8_stage_4_0_t73[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t75 = FSM_dct_8x8_stage_4_0_t74 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_4_0_t76 = FSM_dct_8x8_stage_4_0_t75[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t77 = FSM_dct_8x8_stage_4_0_t76[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t78 = i_data_in[FSM_dct_8x8_stage_4_0_t77 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t79 = FSM_dct_8x8_stage_4_0_t78 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t80 = FSM_dct_8x8_stage_4_0_t79[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t81 = FSM_dct_8x8_stage_4_0_t67;
    FSM_dct_8x8_stage_4_0_t81[FSM_dct_8x8_stage_4_0_t72 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t80;
    FSM_dct_8x8_stage_4_0_t82 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_4_0_t83 = FSM_dct_8x8_stage_4_0_t82[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t84 = FSM_dct_8x8_stage_4_0_t83 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_4_0_t85 = FSM_dct_8x8_stage_4_0_t84[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t86 = FSM_dct_8x8_stage_4_0_t85[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t87 = FSM_dct_8x8_stage_4_0_t64 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t88 = FSM_dct_8x8_stage_4_0_t87[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t89 = FSM_dct_8x8_stage_4_0_t81;
    FSM_dct_8x8_stage_4_0_t89[FSM_dct_8x8_stage_4_0_t86 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t88 - FSM_dct_8x8_stage_4_0_t66;
    FSM_dct_8x8_stage_4_0_t90 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_4_0_t91 = FSM_dct_8x8_stage_4_0_t90[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t92 = FSM_dct_8x8_stage_4_0_t91 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_4_0_t93 = FSM_dct_8x8_stage_4_0_t92[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t94 = FSM_dct_8x8_stage_4_0_t93[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t95 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_4_0_t96 = FSM_dct_8x8_stage_4_0_t95[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t97 = FSM_dct_8x8_stage_4_0_t96 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_4_0_t98 = FSM_dct_8x8_stage_4_0_t97[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t99 = FSM_dct_8x8_stage_4_0_t98[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t100 = i_data_in[FSM_dct_8x8_stage_4_0_t99 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t101 = FSM_dct_8x8_stage_4_0_t89;
    FSM_dct_8x8_stage_4_0_t101[FSM_dct_8x8_stage_4_0_t94 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t100;
    FSM_dct_8x8_stage_4_0_t102 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_4_0_t103 = FSM_dct_8x8_stage_4_0_t102[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t104 = FSM_dct_8x8_stage_4_0_t103[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t105 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_4_0_t106 = FSM_dct_8x8_stage_4_0_t105[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t107 = FSM_dct_8x8_stage_4_0_t106[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t108 = i_data_in[FSM_dct_8x8_stage_4_0_t107 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t109 = FSM_dct_8x8_stage_4_0_t101;
    FSM_dct_8x8_stage_4_0_t109[FSM_dct_8x8_stage_4_0_t104 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t108;
    FSM_dct_8x8_stage_4_0_t110 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_4_0_t111 = FSM_dct_8x8_stage_4_0_t110[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t112 = FSM_dct_8x8_stage_4_0_t111 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_4_0_t113 = FSM_dct_8x8_stage_4_0_t112[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t114 = FSM_dct_8x8_stage_4_0_t113[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t115 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_4_0_t116 = FSM_dct_8x8_stage_4_0_t115[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t117 = FSM_dct_8x8_stage_4_0_t116 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_4_0_t118 = FSM_dct_8x8_stage_4_0_t117[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t119 = FSM_dct_8x8_stage_4_0_t118[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t120 = i_data_in[FSM_dct_8x8_stage_4_0_t119 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t121 = FSM_dct_8x8_stage_4_0_t109;
    FSM_dct_8x8_stage_4_0_t121[FSM_dct_8x8_stage_4_0_t114 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t120;
    FSM_dct_8x8_stage_4_0_t122 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_4_0_t123 = FSM_dct_8x8_stage_4_0_t122[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t124 = FSM_dct_8x8_stage_4_0_t123 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_4_0_t125 = FSM_dct_8x8_stage_4_0_t124[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t126 = FSM_dct_8x8_stage_4_0_t125[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t127 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_4_0_t128 = FSM_dct_8x8_stage_4_0_t127[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t129 = FSM_dct_8x8_stage_4_0_t128 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_4_0_t130 = FSM_dct_8x8_stage_4_0_t129[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t131 = FSM_dct_8x8_stage_4_0_t130[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t132 = i_data_in[FSM_dct_8x8_stage_4_0_t131 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t133 = FSM_dct_8x8_stage_4_0_t132 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t134 = FSM_dct_8x8_stage_4_0_t133[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t135 = FSM_dct_8x8_stage_4_0_t121;
    FSM_dct_8x8_stage_4_0_t135[FSM_dct_8x8_stage_4_0_t126 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t134;
    FSM_dct_8x8_stage_4_0_t136 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_4_0_t137 = FSM_dct_8x8_stage_4_0_t136[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t138 = FSM_dct_8x8_stage_4_0_t137 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_4_0_t139 = FSM_dct_8x8_stage_4_0_t138[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t140 = FSM_dct_8x8_stage_4_0_t139[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t141 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_4_0_t142 = FSM_dct_8x8_stage_4_0_t141[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t143 = FSM_dct_8x8_stage_4_0_t142 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_4_0_t144 = FSM_dct_8x8_stage_4_0_t143[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t145 = FSM_dct_8x8_stage_4_0_t144[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t146 = i_data_in[FSM_dct_8x8_stage_4_0_t145 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t147 = FSM_dct_8x8_stage_4_0_t135;
    FSM_dct_8x8_stage_4_0_t147[FSM_dct_8x8_stage_4_0_t140 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t146;
    FSM_dct_8x8_stage_4_0_t148 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_4_0_t149 = FSM_dct_8x8_stage_4_0_t148[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t150 = FSM_dct_8x8_stage_4_0_t149 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_4_0_t151 = FSM_dct_8x8_stage_4_0_t150[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t152 = FSM_dct_8x8_stage_4_0_t151[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t153 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_4_0_t154 = FSM_dct_8x8_stage_4_0_t153[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t155 = FSM_dct_8x8_stage_4_0_t154 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_4_0_t156 = FSM_dct_8x8_stage_4_0_t155[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t157 = FSM_dct_8x8_stage_4_0_t156[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t158 = i_data_in[FSM_dct_8x8_stage_4_0_t157 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t159 = FSM_dct_8x8_stage_4_0_t158 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t160 = FSM_dct_8x8_stage_4_0_t159[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t161 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_4_0_t162 = FSM_dct_8x8_stage_4_0_t161[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t163 = FSM_dct_8x8_stage_4_0_t162 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_4_0_t164 = FSM_dct_8x8_stage_4_0_t163[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t165 = FSM_dct_8x8_stage_4_0_t164[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t166 = i_data_in[FSM_dct_8x8_stage_4_0_t165 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t167 = (FSM_dct_8x8_stage_4_0_t166 - FSM_dct_8x8_stage_4_0_t158) * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t168 = FSM_dct_8x8_stage_4_0_t167[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t169 = FSM_dct_8x8_stage_4_0_t147;
    FSM_dct_8x8_stage_4_0_t169[FSM_dct_8x8_stage_4_0_t152 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t160 - FSM_dct_8x8_stage_4_0_t168;
    FSM_dct_8x8_stage_4_0_t170 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_4_0_t171 = FSM_dct_8x8_stage_4_0_t170[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t172 = FSM_dct_8x8_stage_4_0_t171 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_4_0_t173 = FSM_dct_8x8_stage_4_0_t172[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t174 = FSM_dct_8x8_stage_4_0_t173[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t175 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_4_0_t176 = FSM_dct_8x8_stage_4_0_t175[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t177 = FSM_dct_8x8_stage_4_0_t176 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_4_0_t178 = FSM_dct_8x8_stage_4_0_t177[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t179 = FSM_dct_8x8_stage_4_0_t178[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t180 = i_data_in[FSM_dct_8x8_stage_4_0_t179 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t181 = FSM_dct_8x8_stage_4_0_t180 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t182 = FSM_dct_8x8_stage_4_0_t181[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t183 = FSM_dct_8x8_stage_4_0_t169;
    FSM_dct_8x8_stage_4_0_t183[FSM_dct_8x8_stage_4_0_t174 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t182;
    FSM_dct_8x8_stage_4_0_t184 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_4_0_t185 = FSM_dct_8x8_stage_4_0_t184[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t186 = FSM_dct_8x8_stage_4_0_t185 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_4_0_t187 = FSM_dct_8x8_stage_4_0_t186[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t188 = FSM_dct_8x8_stage_4_0_t187[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t189 = FSM_dct_8x8_stage_4_0_t166 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t190 = FSM_dct_8x8_stage_4_0_t189[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t191 = FSM_dct_8x8_stage_4_0_t183;
    FSM_dct_8x8_stage_4_0_t191[FSM_dct_8x8_stage_4_0_t188 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t190 - FSM_dct_8x8_stage_4_0_t168;
    FSM_dct_8x8_stage_4_0_t192 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_4_0_t193 = FSM_dct_8x8_stage_4_0_t192[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t194 = FSM_dct_8x8_stage_4_0_t193 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_4_0_t195 = FSM_dct_8x8_stage_4_0_t194[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t196 = FSM_dct_8x8_stage_4_0_t195[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t197 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_4_0_t198 = FSM_dct_8x8_stage_4_0_t197[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t199 = FSM_dct_8x8_stage_4_0_t198 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_4_0_t200 = FSM_dct_8x8_stage_4_0_t199[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t201 = FSM_dct_8x8_stage_4_0_t200[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t202 = i_data_in[FSM_dct_8x8_stage_4_0_t201 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t203 = FSM_dct_8x8_stage_4_0_t191;
    FSM_dct_8x8_stage_4_0_t203[FSM_dct_8x8_stage_4_0_t196 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t202;
    FSM_dct_8x8_stage_4_0_t204 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_4_0_t205 = FSM_dct_8x8_stage_4_0_t204[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t206 = FSM_dct_8x8_stage_4_0_t205[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t207 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_4_0_t208 = FSM_dct_8x8_stage_4_0_t207[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t209 = FSM_dct_8x8_stage_4_0_t208[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t210 = i_data_in[FSM_dct_8x8_stage_4_0_t209 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t211 = FSM_dct_8x8_stage_4_0_t203;
    FSM_dct_8x8_stage_4_0_t211[FSM_dct_8x8_stage_4_0_t206 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t210;
    FSM_dct_8x8_stage_4_0_t212 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_4_0_t213 = FSM_dct_8x8_stage_4_0_t212[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t214 = FSM_dct_8x8_stage_4_0_t213 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_4_0_t215 = FSM_dct_8x8_stage_4_0_t214[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t216 = FSM_dct_8x8_stage_4_0_t215[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t217 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_4_0_t218 = FSM_dct_8x8_stage_4_0_t217[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t219 = FSM_dct_8x8_stage_4_0_t218 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_4_0_t220 = FSM_dct_8x8_stage_4_0_t219[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t221 = FSM_dct_8x8_stage_4_0_t220[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t222 = i_data_in[FSM_dct_8x8_stage_4_0_t221 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t223 = FSM_dct_8x8_stage_4_0_t211;
    FSM_dct_8x8_stage_4_0_t223[FSM_dct_8x8_stage_4_0_t216 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t222;
    FSM_dct_8x8_stage_4_0_t224 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_4_0_t225 = FSM_dct_8x8_stage_4_0_t224[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t226 = FSM_dct_8x8_stage_4_0_t225 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_4_0_t227 = FSM_dct_8x8_stage_4_0_t226[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t228 = FSM_dct_8x8_stage_4_0_t227[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t229 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_4_0_t230 = FSM_dct_8x8_stage_4_0_t229[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t231 = FSM_dct_8x8_stage_4_0_t230 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_4_0_t232 = FSM_dct_8x8_stage_4_0_t231[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t233 = FSM_dct_8x8_stage_4_0_t232[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t234 = i_data_in[FSM_dct_8x8_stage_4_0_t233 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t235 = FSM_dct_8x8_stage_4_0_t234 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t236 = FSM_dct_8x8_stage_4_0_t235[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t237 = FSM_dct_8x8_stage_4_0_t223;
    FSM_dct_8x8_stage_4_0_t237[FSM_dct_8x8_stage_4_0_t228 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t236;
    FSM_dct_8x8_stage_4_0_t238 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_4_0_t239 = FSM_dct_8x8_stage_4_0_t238[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t240 = FSM_dct_8x8_stage_4_0_t239 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_4_0_t241 = FSM_dct_8x8_stage_4_0_t240[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t242 = FSM_dct_8x8_stage_4_0_t241[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t243 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_4_0_t244 = FSM_dct_8x8_stage_4_0_t243[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t245 = FSM_dct_8x8_stage_4_0_t244 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_4_0_t246 = FSM_dct_8x8_stage_4_0_t245[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t247 = FSM_dct_8x8_stage_4_0_t246[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t248 = i_data_in[FSM_dct_8x8_stage_4_0_t247 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t249 = FSM_dct_8x8_stage_4_0_t237;
    FSM_dct_8x8_stage_4_0_t249[FSM_dct_8x8_stage_4_0_t242 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t248;
    FSM_dct_8x8_stage_4_0_t250 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_4_0_t251 = FSM_dct_8x8_stage_4_0_t250[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t252 = FSM_dct_8x8_stage_4_0_t251 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_4_0_t253 = FSM_dct_8x8_stage_4_0_t252[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t254 = FSM_dct_8x8_stage_4_0_t253[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t255 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_4_0_t256 = FSM_dct_8x8_stage_4_0_t255[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t257 = FSM_dct_8x8_stage_4_0_t256 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_4_0_t258 = FSM_dct_8x8_stage_4_0_t257[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t259 = FSM_dct_8x8_stage_4_0_t258[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t260 = i_data_in[FSM_dct_8x8_stage_4_0_t259 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t261 = FSM_dct_8x8_stage_4_0_t260 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t262 = FSM_dct_8x8_stage_4_0_t261[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t263 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_4_0_t264 = FSM_dct_8x8_stage_4_0_t263[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t265 = FSM_dct_8x8_stage_4_0_t264 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_4_0_t266 = FSM_dct_8x8_stage_4_0_t265[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t267 = FSM_dct_8x8_stage_4_0_t266[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t268 = i_data_in[FSM_dct_8x8_stage_4_0_t267 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t269 = (FSM_dct_8x8_stage_4_0_t268 - FSM_dct_8x8_stage_4_0_t260) * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t270 = FSM_dct_8x8_stage_4_0_t269[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t271 = FSM_dct_8x8_stage_4_0_t249;
    FSM_dct_8x8_stage_4_0_t271[FSM_dct_8x8_stage_4_0_t254 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t262 - FSM_dct_8x8_stage_4_0_t270;
    FSM_dct_8x8_stage_4_0_t272 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_4_0_t273 = FSM_dct_8x8_stage_4_0_t272[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t274 = FSM_dct_8x8_stage_4_0_t273 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_4_0_t275 = FSM_dct_8x8_stage_4_0_t274[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t276 = FSM_dct_8x8_stage_4_0_t275[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t277 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_4_0_t278 = FSM_dct_8x8_stage_4_0_t277[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t279 = FSM_dct_8x8_stage_4_0_t278 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_4_0_t280 = FSM_dct_8x8_stage_4_0_t279[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t281 = FSM_dct_8x8_stage_4_0_t280[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t282 = i_data_in[FSM_dct_8x8_stage_4_0_t281 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t283 = FSM_dct_8x8_stage_4_0_t282 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t284 = FSM_dct_8x8_stage_4_0_t283[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t285 = FSM_dct_8x8_stage_4_0_t271;
    FSM_dct_8x8_stage_4_0_t285[FSM_dct_8x8_stage_4_0_t276 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t284;
    FSM_dct_8x8_stage_4_0_t286 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_4_0_t287 = FSM_dct_8x8_stage_4_0_t286[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t288 = FSM_dct_8x8_stage_4_0_t287 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_4_0_t289 = FSM_dct_8x8_stage_4_0_t288[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t290 = FSM_dct_8x8_stage_4_0_t289[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t291 = FSM_dct_8x8_stage_4_0_t268 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t292 = FSM_dct_8x8_stage_4_0_t291[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t293 = FSM_dct_8x8_stage_4_0_t285;
    FSM_dct_8x8_stage_4_0_t293[FSM_dct_8x8_stage_4_0_t290 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t292 - FSM_dct_8x8_stage_4_0_t270;
    FSM_dct_8x8_stage_4_0_t294 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_4_0_t295 = FSM_dct_8x8_stage_4_0_t294[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t296 = FSM_dct_8x8_stage_4_0_t295 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_4_0_t297 = FSM_dct_8x8_stage_4_0_t296[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t298 = FSM_dct_8x8_stage_4_0_t297[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t299 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_4_0_t300 = FSM_dct_8x8_stage_4_0_t299[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t301 = FSM_dct_8x8_stage_4_0_t300 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_4_0_t302 = FSM_dct_8x8_stage_4_0_t301[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t303 = FSM_dct_8x8_stage_4_0_t302[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t304 = i_data_in[FSM_dct_8x8_stage_4_0_t303 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t305 = FSM_dct_8x8_stage_4_0_t293;
    FSM_dct_8x8_stage_4_0_t305[FSM_dct_8x8_stage_4_0_t298 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t304;
    FSM_dct_8x8_stage_4_0_t306 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_4_0_t307 = FSM_dct_8x8_stage_4_0_t306[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t308 = FSM_dct_8x8_stage_4_0_t307[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t309 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_4_0_t310 = FSM_dct_8x8_stage_4_0_t309[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t311 = FSM_dct_8x8_stage_4_0_t310[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t312 = i_data_in[FSM_dct_8x8_stage_4_0_t311 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t313 = FSM_dct_8x8_stage_4_0_t305;
    FSM_dct_8x8_stage_4_0_t313[FSM_dct_8x8_stage_4_0_t308 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t312;
    FSM_dct_8x8_stage_4_0_t314 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_4_0_t315 = FSM_dct_8x8_stage_4_0_t314[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t316 = FSM_dct_8x8_stage_4_0_t315 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_4_0_t317 = FSM_dct_8x8_stage_4_0_t316[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t318 = FSM_dct_8x8_stage_4_0_t317[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t319 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_4_0_t320 = FSM_dct_8x8_stage_4_0_t319[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t321 = FSM_dct_8x8_stage_4_0_t320 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_4_0_t322 = FSM_dct_8x8_stage_4_0_t321[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t323 = FSM_dct_8x8_stage_4_0_t322[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t324 = i_data_in[FSM_dct_8x8_stage_4_0_t323 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t325 = FSM_dct_8x8_stage_4_0_t313;
    FSM_dct_8x8_stage_4_0_t325[FSM_dct_8x8_stage_4_0_t318 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t324;
    FSM_dct_8x8_stage_4_0_t326 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_4_0_t327 = FSM_dct_8x8_stage_4_0_t326[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t328 = FSM_dct_8x8_stage_4_0_t327 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_4_0_t329 = FSM_dct_8x8_stage_4_0_t328[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t330 = FSM_dct_8x8_stage_4_0_t329[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t331 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_4_0_t332 = FSM_dct_8x8_stage_4_0_t331[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t333 = FSM_dct_8x8_stage_4_0_t332 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_4_0_t334 = FSM_dct_8x8_stage_4_0_t333[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t335 = FSM_dct_8x8_stage_4_0_t334[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t336 = i_data_in[FSM_dct_8x8_stage_4_0_t335 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t337 = FSM_dct_8x8_stage_4_0_t336 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t338 = FSM_dct_8x8_stage_4_0_t337[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t339 = FSM_dct_8x8_stage_4_0_t325;
    FSM_dct_8x8_stage_4_0_t339[FSM_dct_8x8_stage_4_0_t330 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t338;
    FSM_dct_8x8_stage_4_0_t340 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_4_0_t341 = FSM_dct_8x8_stage_4_0_t340[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t342 = FSM_dct_8x8_stage_4_0_t341 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_4_0_t343 = FSM_dct_8x8_stage_4_0_t342[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t344 = FSM_dct_8x8_stage_4_0_t343[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t345 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_4_0_t346 = FSM_dct_8x8_stage_4_0_t345[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t347 = FSM_dct_8x8_stage_4_0_t346 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_4_0_t348 = FSM_dct_8x8_stage_4_0_t347[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t349 = FSM_dct_8x8_stage_4_0_t348[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t350 = i_data_in[FSM_dct_8x8_stage_4_0_t349 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t351 = FSM_dct_8x8_stage_4_0_t339;
    FSM_dct_8x8_stage_4_0_t351[FSM_dct_8x8_stage_4_0_t344 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t350;
    FSM_dct_8x8_stage_4_0_t352 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_4_0_t353 = FSM_dct_8x8_stage_4_0_t352[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t354 = FSM_dct_8x8_stage_4_0_t353 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_4_0_t355 = FSM_dct_8x8_stage_4_0_t354[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t356 = FSM_dct_8x8_stage_4_0_t355[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t357 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_4_0_t358 = FSM_dct_8x8_stage_4_0_t357[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t359 = FSM_dct_8x8_stage_4_0_t358 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_4_0_t360 = FSM_dct_8x8_stage_4_0_t359[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t361 = FSM_dct_8x8_stage_4_0_t360[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t362 = i_data_in[FSM_dct_8x8_stage_4_0_t361 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t363 = FSM_dct_8x8_stage_4_0_t362 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t364 = FSM_dct_8x8_stage_4_0_t363[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t365 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_4_0_t366 = FSM_dct_8x8_stage_4_0_t365[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t367 = FSM_dct_8x8_stage_4_0_t366 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_4_0_t368 = FSM_dct_8x8_stage_4_0_t367[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t369 = FSM_dct_8x8_stage_4_0_t368[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t370 = i_data_in[FSM_dct_8x8_stage_4_0_t369 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t371 = (FSM_dct_8x8_stage_4_0_t370 - FSM_dct_8x8_stage_4_0_t362) * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t372 = FSM_dct_8x8_stage_4_0_t371[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t373 = FSM_dct_8x8_stage_4_0_t351;
    FSM_dct_8x8_stage_4_0_t373[FSM_dct_8x8_stage_4_0_t356 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t364 - FSM_dct_8x8_stage_4_0_t372;
    FSM_dct_8x8_stage_4_0_t374 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_4_0_t375 = FSM_dct_8x8_stage_4_0_t374[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t376 = FSM_dct_8x8_stage_4_0_t375 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_4_0_t377 = FSM_dct_8x8_stage_4_0_t376[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t378 = FSM_dct_8x8_stage_4_0_t377[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t379 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_4_0_t380 = FSM_dct_8x8_stage_4_0_t379[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t381 = FSM_dct_8x8_stage_4_0_t380 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_4_0_t382 = FSM_dct_8x8_stage_4_0_t381[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t383 = FSM_dct_8x8_stage_4_0_t382[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t384 = i_data_in[FSM_dct_8x8_stage_4_0_t383 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t385 = FSM_dct_8x8_stage_4_0_t384 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t386 = FSM_dct_8x8_stage_4_0_t385[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t387 = FSM_dct_8x8_stage_4_0_t373;
    FSM_dct_8x8_stage_4_0_t387[FSM_dct_8x8_stage_4_0_t378 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t386;
    FSM_dct_8x8_stage_4_0_t388 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_4_0_t389 = FSM_dct_8x8_stage_4_0_t388[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t390 = FSM_dct_8x8_stage_4_0_t389 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_4_0_t391 = FSM_dct_8x8_stage_4_0_t390[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t392 = FSM_dct_8x8_stage_4_0_t391[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t393 = FSM_dct_8x8_stage_4_0_t370 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t394 = FSM_dct_8x8_stage_4_0_t393[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t395 = FSM_dct_8x8_stage_4_0_t387;
    FSM_dct_8x8_stage_4_0_t395[FSM_dct_8x8_stage_4_0_t392 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t394 - FSM_dct_8x8_stage_4_0_t372;
    FSM_dct_8x8_stage_4_0_t396 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_4_0_t397 = FSM_dct_8x8_stage_4_0_t396[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t398 = FSM_dct_8x8_stage_4_0_t397 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_4_0_t399 = FSM_dct_8x8_stage_4_0_t398[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t400 = FSM_dct_8x8_stage_4_0_t399[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t401 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_4_0_t402 = FSM_dct_8x8_stage_4_0_t401[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t403 = FSM_dct_8x8_stage_4_0_t402 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_4_0_t404 = FSM_dct_8x8_stage_4_0_t403[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t405 = FSM_dct_8x8_stage_4_0_t404[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t406 = i_data_in[FSM_dct_8x8_stage_4_0_t405 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t407 = FSM_dct_8x8_stage_4_0_t395;
    FSM_dct_8x8_stage_4_0_t407[FSM_dct_8x8_stage_4_0_t400 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t406;
    FSM_dct_8x8_stage_4_0_t408 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_4_0_t409 = FSM_dct_8x8_stage_4_0_t408[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t410 = FSM_dct_8x8_stage_4_0_t409[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t411 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_4_0_t412 = FSM_dct_8x8_stage_4_0_t411[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t413 = FSM_dct_8x8_stage_4_0_t412[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t414 = i_data_in[FSM_dct_8x8_stage_4_0_t413 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t415 = FSM_dct_8x8_stage_4_0_t407;
    FSM_dct_8x8_stage_4_0_t415[FSM_dct_8x8_stage_4_0_t410 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t414;
    FSM_dct_8x8_stage_4_0_t416 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_4_0_t417 = FSM_dct_8x8_stage_4_0_t416[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t418 = FSM_dct_8x8_stage_4_0_t417 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_4_0_t419 = FSM_dct_8x8_stage_4_0_t418[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t420 = FSM_dct_8x8_stage_4_0_t419[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t421 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_4_0_t422 = FSM_dct_8x8_stage_4_0_t421[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t423 = FSM_dct_8x8_stage_4_0_t422 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_4_0_t424 = FSM_dct_8x8_stage_4_0_t423[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t425 = FSM_dct_8x8_stage_4_0_t424[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t426 = i_data_in[FSM_dct_8x8_stage_4_0_t425 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t427 = FSM_dct_8x8_stage_4_0_t415;
    FSM_dct_8x8_stage_4_0_t427[FSM_dct_8x8_stage_4_0_t420 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t426;
    FSM_dct_8x8_stage_4_0_t428 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_4_0_t429 = FSM_dct_8x8_stage_4_0_t428[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t430 = FSM_dct_8x8_stage_4_0_t429 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_4_0_t431 = FSM_dct_8x8_stage_4_0_t430[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t432 = FSM_dct_8x8_stage_4_0_t431[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t433 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_4_0_t434 = FSM_dct_8x8_stage_4_0_t433[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t435 = FSM_dct_8x8_stage_4_0_t434 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_4_0_t436 = FSM_dct_8x8_stage_4_0_t435[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t437 = FSM_dct_8x8_stage_4_0_t436[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t438 = i_data_in[FSM_dct_8x8_stage_4_0_t437 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t439 = FSM_dct_8x8_stage_4_0_t438 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t440 = FSM_dct_8x8_stage_4_0_t439[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t441 = FSM_dct_8x8_stage_4_0_t427;
    FSM_dct_8x8_stage_4_0_t441[FSM_dct_8x8_stage_4_0_t432 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t440;
    FSM_dct_8x8_stage_4_0_t442 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_4_0_t443 = FSM_dct_8x8_stage_4_0_t442[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t444 = FSM_dct_8x8_stage_4_0_t443 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_4_0_t445 = FSM_dct_8x8_stage_4_0_t444[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t446 = FSM_dct_8x8_stage_4_0_t445[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t447 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_4_0_t448 = FSM_dct_8x8_stage_4_0_t447[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t449 = FSM_dct_8x8_stage_4_0_t448 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_4_0_t450 = FSM_dct_8x8_stage_4_0_t449[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t451 = FSM_dct_8x8_stage_4_0_t450[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t452 = i_data_in[FSM_dct_8x8_stage_4_0_t451 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t453 = FSM_dct_8x8_stage_4_0_t441;
    FSM_dct_8x8_stage_4_0_t453[FSM_dct_8x8_stage_4_0_t446 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t452;
    FSM_dct_8x8_stage_4_0_t454 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_4_0_t455 = FSM_dct_8x8_stage_4_0_t454[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t456 = FSM_dct_8x8_stage_4_0_t455 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_4_0_t457 = FSM_dct_8x8_stage_4_0_t456[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t458 = FSM_dct_8x8_stage_4_0_t457[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t459 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_4_0_t460 = FSM_dct_8x8_stage_4_0_t459[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t461 = FSM_dct_8x8_stage_4_0_t460 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_4_0_t462 = FSM_dct_8x8_stage_4_0_t461[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t463 = FSM_dct_8x8_stage_4_0_t462[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t464 = i_data_in[FSM_dct_8x8_stage_4_0_t463 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t465 = FSM_dct_8x8_stage_4_0_t464 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t466 = FSM_dct_8x8_stage_4_0_t465[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t467 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_4_0_t468 = FSM_dct_8x8_stage_4_0_t467[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t469 = FSM_dct_8x8_stage_4_0_t468 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_4_0_t470 = FSM_dct_8x8_stage_4_0_t469[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t471 = FSM_dct_8x8_stage_4_0_t470[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t472 = i_data_in[FSM_dct_8x8_stage_4_0_t471 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t473 = (FSM_dct_8x8_stage_4_0_t472 - FSM_dct_8x8_stage_4_0_t464) * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t474 = FSM_dct_8x8_stage_4_0_t473[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t475 = FSM_dct_8x8_stage_4_0_t453;
    FSM_dct_8x8_stage_4_0_t475[FSM_dct_8x8_stage_4_0_t458 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t466 - FSM_dct_8x8_stage_4_0_t474;
    FSM_dct_8x8_stage_4_0_t476 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_4_0_t477 = FSM_dct_8x8_stage_4_0_t476[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t478 = FSM_dct_8x8_stage_4_0_t477 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_4_0_t479 = FSM_dct_8x8_stage_4_0_t478[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t480 = FSM_dct_8x8_stage_4_0_t479[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t481 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_4_0_t482 = FSM_dct_8x8_stage_4_0_t481[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t483 = FSM_dct_8x8_stage_4_0_t482 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_4_0_t484 = FSM_dct_8x8_stage_4_0_t483[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t485 = FSM_dct_8x8_stage_4_0_t484[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t486 = i_data_in[FSM_dct_8x8_stage_4_0_t485 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t487 = FSM_dct_8x8_stage_4_0_t486 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t488 = FSM_dct_8x8_stage_4_0_t487[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t489 = FSM_dct_8x8_stage_4_0_t475;
    FSM_dct_8x8_stage_4_0_t489[FSM_dct_8x8_stage_4_0_t480 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t488;
    FSM_dct_8x8_stage_4_0_t490 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_4_0_t491 = FSM_dct_8x8_stage_4_0_t490[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t492 = FSM_dct_8x8_stage_4_0_t491 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_4_0_t493 = FSM_dct_8x8_stage_4_0_t492[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t494 = FSM_dct_8x8_stage_4_0_t493[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t495 = FSM_dct_8x8_stage_4_0_t472 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t496 = FSM_dct_8x8_stage_4_0_t495[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t497 = FSM_dct_8x8_stage_4_0_t489;
    FSM_dct_8x8_stage_4_0_t497[FSM_dct_8x8_stage_4_0_t494 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t496 - FSM_dct_8x8_stage_4_0_t474;
    FSM_dct_8x8_stage_4_0_t498 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_4_0_t499 = FSM_dct_8x8_stage_4_0_t498[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t500 = FSM_dct_8x8_stage_4_0_t499 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_4_0_t501 = FSM_dct_8x8_stage_4_0_t500[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t502 = FSM_dct_8x8_stage_4_0_t501[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t503 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_4_0_t504 = FSM_dct_8x8_stage_4_0_t503[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t505 = FSM_dct_8x8_stage_4_0_t504 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_4_0_t506 = FSM_dct_8x8_stage_4_0_t505[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t507 = FSM_dct_8x8_stage_4_0_t506[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t508 = i_data_in[FSM_dct_8x8_stage_4_0_t507 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t509 = FSM_dct_8x8_stage_4_0_t497;
    FSM_dct_8x8_stage_4_0_t509[FSM_dct_8x8_stage_4_0_t502 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t508;
    FSM_dct_8x8_stage_4_0_t510 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_4_0_t511 = FSM_dct_8x8_stage_4_0_t510[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t512 = FSM_dct_8x8_stage_4_0_t511[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t513 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_4_0_t514 = FSM_dct_8x8_stage_4_0_t513[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t515 = FSM_dct_8x8_stage_4_0_t514[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t516 = i_data_in[FSM_dct_8x8_stage_4_0_t515 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t517 = FSM_dct_8x8_stage_4_0_t509;
    FSM_dct_8x8_stage_4_0_t517[FSM_dct_8x8_stage_4_0_t512 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t516;
    FSM_dct_8x8_stage_4_0_t518 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_4_0_t519 = FSM_dct_8x8_stage_4_0_t518[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t520 = FSM_dct_8x8_stage_4_0_t519 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_4_0_t521 = FSM_dct_8x8_stage_4_0_t520[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t522 = FSM_dct_8x8_stage_4_0_t521[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t523 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_4_0_t524 = FSM_dct_8x8_stage_4_0_t523[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t525 = FSM_dct_8x8_stage_4_0_t524 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_4_0_t526 = FSM_dct_8x8_stage_4_0_t525[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t527 = FSM_dct_8x8_stage_4_0_t526[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t528 = i_data_in[FSM_dct_8x8_stage_4_0_t527 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t529 = FSM_dct_8x8_stage_4_0_t517;
    FSM_dct_8x8_stage_4_0_t529[FSM_dct_8x8_stage_4_0_t522 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t528;
    FSM_dct_8x8_stage_4_0_t530 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_4_0_t531 = FSM_dct_8x8_stage_4_0_t530[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t532 = FSM_dct_8x8_stage_4_0_t531 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_4_0_t533 = FSM_dct_8x8_stage_4_0_t532[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t534 = FSM_dct_8x8_stage_4_0_t533[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t535 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_4_0_t536 = FSM_dct_8x8_stage_4_0_t535[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t537 = FSM_dct_8x8_stage_4_0_t536 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_4_0_t538 = FSM_dct_8x8_stage_4_0_t537[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t539 = FSM_dct_8x8_stage_4_0_t538[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t540 = i_data_in[FSM_dct_8x8_stage_4_0_t539 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t541 = FSM_dct_8x8_stage_4_0_t540 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t542 = FSM_dct_8x8_stage_4_0_t541[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t543 = FSM_dct_8x8_stage_4_0_t529;
    FSM_dct_8x8_stage_4_0_t543[FSM_dct_8x8_stage_4_0_t534 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t542;
    FSM_dct_8x8_stage_4_0_t544 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_4_0_t545 = FSM_dct_8x8_stage_4_0_t544[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t546 = FSM_dct_8x8_stage_4_0_t545 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_4_0_t547 = FSM_dct_8x8_stage_4_0_t546[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t548 = FSM_dct_8x8_stage_4_0_t547[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t549 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_4_0_t550 = FSM_dct_8x8_stage_4_0_t549[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t551 = FSM_dct_8x8_stage_4_0_t550 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_4_0_t552 = FSM_dct_8x8_stage_4_0_t551[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t553 = FSM_dct_8x8_stage_4_0_t552[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t554 = i_data_in[FSM_dct_8x8_stage_4_0_t553 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t555 = FSM_dct_8x8_stage_4_0_t543;
    FSM_dct_8x8_stage_4_0_t555[FSM_dct_8x8_stage_4_0_t548 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t554;
    FSM_dct_8x8_stage_4_0_t556 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_4_0_t557 = FSM_dct_8x8_stage_4_0_t556[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t558 = FSM_dct_8x8_stage_4_0_t557 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_4_0_t559 = FSM_dct_8x8_stage_4_0_t558[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t560 = FSM_dct_8x8_stage_4_0_t559[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t561 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_4_0_t562 = FSM_dct_8x8_stage_4_0_t561[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t563 = FSM_dct_8x8_stage_4_0_t562 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_4_0_t564 = FSM_dct_8x8_stage_4_0_t563[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t565 = FSM_dct_8x8_stage_4_0_t564[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t566 = i_data_in[FSM_dct_8x8_stage_4_0_t565 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t567 = FSM_dct_8x8_stage_4_0_t566 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t568 = FSM_dct_8x8_stage_4_0_t567[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t569 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_4_0_t570 = FSM_dct_8x8_stage_4_0_t569[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t571 = FSM_dct_8x8_stage_4_0_t570 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_4_0_t572 = FSM_dct_8x8_stage_4_0_t571[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t573 = FSM_dct_8x8_stage_4_0_t572[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t574 = i_data_in[FSM_dct_8x8_stage_4_0_t573 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t575 = (FSM_dct_8x8_stage_4_0_t574 - FSM_dct_8x8_stage_4_0_t566) * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t576 = FSM_dct_8x8_stage_4_0_t575[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t577 = FSM_dct_8x8_stage_4_0_t555;
    FSM_dct_8x8_stage_4_0_t577[FSM_dct_8x8_stage_4_0_t560 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t568 - FSM_dct_8x8_stage_4_0_t576;
    FSM_dct_8x8_stage_4_0_t578 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_4_0_t579 = FSM_dct_8x8_stage_4_0_t578[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t580 = FSM_dct_8x8_stage_4_0_t579 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_4_0_t581 = FSM_dct_8x8_stage_4_0_t580[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t582 = FSM_dct_8x8_stage_4_0_t581[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t583 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_4_0_t584 = FSM_dct_8x8_stage_4_0_t583[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t585 = FSM_dct_8x8_stage_4_0_t584 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_4_0_t586 = FSM_dct_8x8_stage_4_0_t585[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t587 = FSM_dct_8x8_stage_4_0_t586[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t588 = i_data_in[FSM_dct_8x8_stage_4_0_t587 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t589 = FSM_dct_8x8_stage_4_0_t588 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t590 = FSM_dct_8x8_stage_4_0_t589[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t591 = FSM_dct_8x8_stage_4_0_t577;
    FSM_dct_8x8_stage_4_0_t591[FSM_dct_8x8_stage_4_0_t582 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t590;
    FSM_dct_8x8_stage_4_0_t592 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_4_0_t593 = FSM_dct_8x8_stage_4_0_t592[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t594 = FSM_dct_8x8_stage_4_0_t593 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_4_0_t595 = FSM_dct_8x8_stage_4_0_t594[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t596 = FSM_dct_8x8_stage_4_0_t595[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t597 = FSM_dct_8x8_stage_4_0_t574 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t598 = FSM_dct_8x8_stage_4_0_t597[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t599 = FSM_dct_8x8_stage_4_0_t591;
    FSM_dct_8x8_stage_4_0_t599[FSM_dct_8x8_stage_4_0_t596 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t598 - FSM_dct_8x8_stage_4_0_t576;
    FSM_dct_8x8_stage_4_0_t600 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_4_0_t601 = FSM_dct_8x8_stage_4_0_t600[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t602 = FSM_dct_8x8_stage_4_0_t601 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_4_0_t603 = FSM_dct_8x8_stage_4_0_t602[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t604 = FSM_dct_8x8_stage_4_0_t603[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t605 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_4_0_t606 = FSM_dct_8x8_stage_4_0_t605[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t607 = FSM_dct_8x8_stage_4_0_t606 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_4_0_t608 = FSM_dct_8x8_stage_4_0_t607[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t609 = FSM_dct_8x8_stage_4_0_t608[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t610 = i_data_in[FSM_dct_8x8_stage_4_0_t609 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t611 = FSM_dct_8x8_stage_4_0_t599;
    FSM_dct_8x8_stage_4_0_t611[FSM_dct_8x8_stage_4_0_t604 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t610;
    FSM_dct_8x8_stage_4_0_t612 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_4_0_t613 = FSM_dct_8x8_stage_4_0_t612[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t614 = FSM_dct_8x8_stage_4_0_t613[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t615 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_4_0_t616 = FSM_dct_8x8_stage_4_0_t615[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t617 = FSM_dct_8x8_stage_4_0_t616[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t618 = i_data_in[FSM_dct_8x8_stage_4_0_t617 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t619 = FSM_dct_8x8_stage_4_0_t611;
    FSM_dct_8x8_stage_4_0_t619[FSM_dct_8x8_stage_4_0_t614 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t618;
    FSM_dct_8x8_stage_4_0_t620 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_4_0_t621 = FSM_dct_8x8_stage_4_0_t620[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t622 = FSM_dct_8x8_stage_4_0_t621 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_4_0_t623 = FSM_dct_8x8_stage_4_0_t622[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t624 = FSM_dct_8x8_stage_4_0_t623[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t625 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_4_0_t626 = FSM_dct_8x8_stage_4_0_t625[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t627 = FSM_dct_8x8_stage_4_0_t626 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_4_0_t628 = FSM_dct_8x8_stage_4_0_t627[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t629 = FSM_dct_8x8_stage_4_0_t628[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t630 = i_data_in[FSM_dct_8x8_stage_4_0_t629 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t631 = FSM_dct_8x8_stage_4_0_t619;
    FSM_dct_8x8_stage_4_0_t631[FSM_dct_8x8_stage_4_0_t624 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t630;
    FSM_dct_8x8_stage_4_0_t632 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_4_0_t633 = FSM_dct_8x8_stage_4_0_t632[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t634 = FSM_dct_8x8_stage_4_0_t633 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_4_0_t635 = FSM_dct_8x8_stage_4_0_t634[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t636 = FSM_dct_8x8_stage_4_0_t635[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t637 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_4_0_t638 = FSM_dct_8x8_stage_4_0_t637[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t639 = FSM_dct_8x8_stage_4_0_t638 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_4_0_t640 = FSM_dct_8x8_stage_4_0_t639[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t641 = FSM_dct_8x8_stage_4_0_t640[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t642 = i_data_in[FSM_dct_8x8_stage_4_0_t641 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t643 = FSM_dct_8x8_stage_4_0_t642 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t644 = FSM_dct_8x8_stage_4_0_t643[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t645 = FSM_dct_8x8_stage_4_0_t631;
    FSM_dct_8x8_stage_4_0_t645[FSM_dct_8x8_stage_4_0_t636 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t644;
    FSM_dct_8x8_stage_4_0_t646 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_4_0_t647 = FSM_dct_8x8_stage_4_0_t646[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t648 = FSM_dct_8x8_stage_4_0_t647 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_4_0_t649 = FSM_dct_8x8_stage_4_0_t648[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t650 = FSM_dct_8x8_stage_4_0_t649[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t651 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_4_0_t652 = FSM_dct_8x8_stage_4_0_t651[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t653 = FSM_dct_8x8_stage_4_0_t652 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_4_0_t654 = FSM_dct_8x8_stage_4_0_t653[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t655 = FSM_dct_8x8_stage_4_0_t654[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t656 = i_data_in[FSM_dct_8x8_stage_4_0_t655 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t657 = FSM_dct_8x8_stage_4_0_t645;
    FSM_dct_8x8_stage_4_0_t657[FSM_dct_8x8_stage_4_0_t650 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t656;
    FSM_dct_8x8_stage_4_0_t658 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_4_0_t659 = FSM_dct_8x8_stage_4_0_t658[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t660 = FSM_dct_8x8_stage_4_0_t659 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_4_0_t661 = FSM_dct_8x8_stage_4_0_t660[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t662 = FSM_dct_8x8_stage_4_0_t661[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t663 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_4_0_t664 = FSM_dct_8x8_stage_4_0_t663[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t665 = FSM_dct_8x8_stage_4_0_t664 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_4_0_t666 = FSM_dct_8x8_stage_4_0_t665[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t667 = FSM_dct_8x8_stage_4_0_t666[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t668 = i_data_in[FSM_dct_8x8_stage_4_0_t667 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t669 = FSM_dct_8x8_stage_4_0_t668 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t670 = FSM_dct_8x8_stage_4_0_t669[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t671 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_4_0_t672 = FSM_dct_8x8_stage_4_0_t671[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t673 = FSM_dct_8x8_stage_4_0_t672 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_4_0_t674 = FSM_dct_8x8_stage_4_0_t673[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t675 = FSM_dct_8x8_stage_4_0_t674[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t676 = i_data_in[FSM_dct_8x8_stage_4_0_t675 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t677 = (FSM_dct_8x8_stage_4_0_t676 - FSM_dct_8x8_stage_4_0_t668) * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t678 = FSM_dct_8x8_stage_4_0_t677[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t679 = FSM_dct_8x8_stage_4_0_t657;
    FSM_dct_8x8_stage_4_0_t679[FSM_dct_8x8_stage_4_0_t662 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t670 - FSM_dct_8x8_stage_4_0_t678;
    FSM_dct_8x8_stage_4_0_t680 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_4_0_t681 = FSM_dct_8x8_stage_4_0_t680[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t682 = FSM_dct_8x8_stage_4_0_t681 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_4_0_t683 = FSM_dct_8x8_stage_4_0_t682[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t684 = FSM_dct_8x8_stage_4_0_t683[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t685 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_4_0_t686 = FSM_dct_8x8_stage_4_0_t685[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t687 = FSM_dct_8x8_stage_4_0_t686 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_4_0_t688 = FSM_dct_8x8_stage_4_0_t687[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t689 = FSM_dct_8x8_stage_4_0_t688[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t690 = i_data_in[FSM_dct_8x8_stage_4_0_t689 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t691 = FSM_dct_8x8_stage_4_0_t690 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t692 = FSM_dct_8x8_stage_4_0_t691[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t693 = FSM_dct_8x8_stage_4_0_t679;
    FSM_dct_8x8_stage_4_0_t693[FSM_dct_8x8_stage_4_0_t684 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t692;
    FSM_dct_8x8_stage_4_0_t694 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_4_0_t695 = FSM_dct_8x8_stage_4_0_t694[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t696 = FSM_dct_8x8_stage_4_0_t695 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_4_0_t697 = FSM_dct_8x8_stage_4_0_t696[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t698 = FSM_dct_8x8_stage_4_0_t697[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t699 = FSM_dct_8x8_stage_4_0_t676 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t700 = FSM_dct_8x8_stage_4_0_t699[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t701 = FSM_dct_8x8_stage_4_0_t693;
    FSM_dct_8x8_stage_4_0_t701[FSM_dct_8x8_stage_4_0_t698 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t700 - FSM_dct_8x8_stage_4_0_t678;
    FSM_dct_8x8_stage_4_0_t702 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_4_0_t703 = FSM_dct_8x8_stage_4_0_t702[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t704 = FSM_dct_8x8_stage_4_0_t703 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_4_0_t705 = FSM_dct_8x8_stage_4_0_t704[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t706 = FSM_dct_8x8_stage_4_0_t705[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t707 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_4_0_t708 = FSM_dct_8x8_stage_4_0_t707[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t709 = FSM_dct_8x8_stage_4_0_t708 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_4_0_t710 = FSM_dct_8x8_stage_4_0_t709[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t711 = FSM_dct_8x8_stage_4_0_t710[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t712 = i_data_in[FSM_dct_8x8_stage_4_0_t711 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t713 = FSM_dct_8x8_stage_4_0_t701;
    FSM_dct_8x8_stage_4_0_t713[FSM_dct_8x8_stage_4_0_t706 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t712;
    FSM_dct_8x8_stage_4_0_t714 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_4_0_t715 = FSM_dct_8x8_stage_4_0_t714[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t716 = FSM_dct_8x8_stage_4_0_t715[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t717 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_4_0_t718 = FSM_dct_8x8_stage_4_0_t717[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t719 = FSM_dct_8x8_stage_4_0_t718[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t720 = i_data_in[FSM_dct_8x8_stage_4_0_t719 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t721 = FSM_dct_8x8_stage_4_0_t713;
    FSM_dct_8x8_stage_4_0_t721[FSM_dct_8x8_stage_4_0_t716 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t720;
    FSM_dct_8x8_stage_4_0_t722 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_4_0_t723 = FSM_dct_8x8_stage_4_0_t722[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t724 = FSM_dct_8x8_stage_4_0_t723 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_4_0_t725 = FSM_dct_8x8_stage_4_0_t724[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t726 = FSM_dct_8x8_stage_4_0_t725[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t727 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_4_0_t728 = FSM_dct_8x8_stage_4_0_t727[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t729 = FSM_dct_8x8_stage_4_0_t728 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_4_0_t730 = FSM_dct_8x8_stage_4_0_t729[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t731 = FSM_dct_8x8_stage_4_0_t730[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t732 = i_data_in[FSM_dct_8x8_stage_4_0_t731 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t733 = FSM_dct_8x8_stage_4_0_t721;
    FSM_dct_8x8_stage_4_0_t733[FSM_dct_8x8_stage_4_0_t726 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t732;
    FSM_dct_8x8_stage_4_0_t734 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_4_0_t735 = FSM_dct_8x8_stage_4_0_t734[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t736 = FSM_dct_8x8_stage_4_0_t735 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_4_0_t737 = FSM_dct_8x8_stage_4_0_t736[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t738 = FSM_dct_8x8_stage_4_0_t737[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t739 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_4_0_t740 = FSM_dct_8x8_stage_4_0_t739[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t741 = FSM_dct_8x8_stage_4_0_t740 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_4_0_t742 = FSM_dct_8x8_stage_4_0_t741[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t743 = FSM_dct_8x8_stage_4_0_t742[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t744 = i_data_in[FSM_dct_8x8_stage_4_0_t743 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t745 = FSM_dct_8x8_stage_4_0_t744 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t746 = FSM_dct_8x8_stage_4_0_t745[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t747 = FSM_dct_8x8_stage_4_0_t733;
    FSM_dct_8x8_stage_4_0_t747[FSM_dct_8x8_stage_4_0_t738 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t746;
    FSM_dct_8x8_stage_4_0_t748 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_4_0_t749 = FSM_dct_8x8_stage_4_0_t748[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t750 = FSM_dct_8x8_stage_4_0_t749 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_4_0_t751 = FSM_dct_8x8_stage_4_0_t750[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t752 = FSM_dct_8x8_stage_4_0_t751[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t753 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_4_0_t754 = FSM_dct_8x8_stage_4_0_t753[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t755 = FSM_dct_8x8_stage_4_0_t754 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_4_0_t756 = FSM_dct_8x8_stage_4_0_t755[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t757 = FSM_dct_8x8_stage_4_0_t756[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t758 = i_data_in[FSM_dct_8x8_stage_4_0_t757 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t759 = FSM_dct_8x8_stage_4_0_t747;
    FSM_dct_8x8_stage_4_0_t759[FSM_dct_8x8_stage_4_0_t752 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t758;
    FSM_dct_8x8_stage_4_0_t760 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_4_0_t761 = FSM_dct_8x8_stage_4_0_t760[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t762 = FSM_dct_8x8_stage_4_0_t761 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_4_0_t763 = FSM_dct_8x8_stage_4_0_t762[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t764 = FSM_dct_8x8_stage_4_0_t763[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t765 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_4_0_t766 = FSM_dct_8x8_stage_4_0_t765[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t767 = FSM_dct_8x8_stage_4_0_t766 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_4_0_t768 = FSM_dct_8x8_stage_4_0_t767[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t769 = FSM_dct_8x8_stage_4_0_t768[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t770 = i_data_in[FSM_dct_8x8_stage_4_0_t769 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t771 = FSM_dct_8x8_stage_4_0_t770 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t772 = FSM_dct_8x8_stage_4_0_t771[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t773 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_4_0_t774 = FSM_dct_8x8_stage_4_0_t773[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t775 = FSM_dct_8x8_stage_4_0_t774 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_4_0_t776 = FSM_dct_8x8_stage_4_0_t775[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t777 = FSM_dct_8x8_stage_4_0_t776[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t778 = i_data_in[FSM_dct_8x8_stage_4_0_t777 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t779 = (FSM_dct_8x8_stage_4_0_t778 - FSM_dct_8x8_stage_4_0_t770) * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t780 = FSM_dct_8x8_stage_4_0_t779[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t781 = FSM_dct_8x8_stage_4_0_t759;
    FSM_dct_8x8_stage_4_0_t781[FSM_dct_8x8_stage_4_0_t764 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t772 - FSM_dct_8x8_stage_4_0_t780;
    FSM_dct_8x8_stage_4_0_t782 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_4_0_t783 = FSM_dct_8x8_stage_4_0_t782[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t784 = FSM_dct_8x8_stage_4_0_t783 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_4_0_t785 = FSM_dct_8x8_stage_4_0_t784[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t786 = FSM_dct_8x8_stage_4_0_t785[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t787 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_4_0_t788 = FSM_dct_8x8_stage_4_0_t787[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t789 = FSM_dct_8x8_stage_4_0_t788 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_4_0_t790 = FSM_dct_8x8_stage_4_0_t789[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t791 = FSM_dct_8x8_stage_4_0_t790[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t792 = i_data_in[FSM_dct_8x8_stage_4_0_t791 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t793 = FSM_dct_8x8_stage_4_0_t792 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t794 = FSM_dct_8x8_stage_4_0_t793[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t795 = FSM_dct_8x8_stage_4_0_t781;
    FSM_dct_8x8_stage_4_0_t795[FSM_dct_8x8_stage_4_0_t786 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t794;
    FSM_dct_8x8_stage_4_0_t796 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_4_0_t797 = FSM_dct_8x8_stage_4_0_t796[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t798 = FSM_dct_8x8_stage_4_0_t797 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_4_0_t799 = FSM_dct_8x8_stage_4_0_t798[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t800 = FSM_dct_8x8_stage_4_0_t799[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t801 = FSM_dct_8x8_stage_4_0_t778 * 32'b00000000000000000000000000010000;
    FSM_dct_8x8_stage_4_0_t802 = FSM_dct_8x8_stage_4_0_t801[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t803 = FSM_dct_8x8_stage_4_0_t795;
    FSM_dct_8x8_stage_4_0_t803[FSM_dct_8x8_stage_4_0_t800 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t802 - FSM_dct_8x8_stage_4_0_t780;
    FSM_dct_8x8_stage_4_0_t804 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_4_0_t805 = FSM_dct_8x8_stage_4_0_t804[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t806 = FSM_dct_8x8_stage_4_0_t805 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_4_0_t807 = FSM_dct_8x8_stage_4_0_t806[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t808 = FSM_dct_8x8_stage_4_0_t807[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t809 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_4_0_t810 = FSM_dct_8x8_stage_4_0_t809[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t811 = FSM_dct_8x8_stage_4_0_t810 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_4_0_t812 = FSM_dct_8x8_stage_4_0_t811[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_4_0_t813 = FSM_dct_8x8_stage_4_0_t812[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_4_0_t814 = i_data_in[FSM_dct_8x8_stage_4_0_t813 * 32 +: 32];
    FSM_dct_8x8_stage_4_0_t815 = FSM_dct_8x8_stage_4_0_t803;
    FSM_dct_8x8_stage_4_0_t815[FSM_dct_8x8_stage_4_0_t808 * 32 +: 32] = FSM_dct_8x8_stage_4_0_t814;
end

assign FSM_dct_8x8_stage_4_0_in_ready = 1'b1;

always @(posedge clk) begin
    FSM_dct_8x8_stage_4_0_st_dummy_reg <= FSM_dct_8x8_stage_4_0_st_dummy_reg;
    if (rst) begin
        FSM_dct_8x8_stage_4_0_st_dummy_reg <= 32'b0;
    end
end
/* End submodules of dct_8x8_stage_4 */
/* End module dct_8x8_stage_4 */
endgenerate
endmodule
