`timescale 1ns / 1ps

module dct_8x8_stage_2_inner
(
    input wire clk,
    input wire rst,
    input wire [2048-1:0] i_data_in,
    input wire i_valid,
    output wire i_ready,
    output wire [2048-1:0] o_data_out,
    output wire o_valid,
    input wire o_ready
);

generate
/*
    Begin module dct_8x8_stage_2
*/
/*
    Wires declared by dct_8x8_stage_2
*/
wire FSM_dct_8x8_stage_2_0_in_ready;
wire FSM_dct_8x8_stage_2_0_out_valid;
/* End wires declared by dct_8x8_stage_2 */

/*
    Submodules of dct_8x8_stage_2
*/
reg [32-1:0] FSM_dct_8x8_stage_2_0_st_dummy_reg = 32'b0;

reg [64-1:0] FSM_dct_8x8_stage_2_0_t0;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t1;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t2;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t3;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t4;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t5;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t6;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t7;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t8;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t9;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t10;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t11;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t12;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t13;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t14;
reg [2048-1:0] FSM_dct_8x8_stage_2_0_t15;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t16;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t17;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t18;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t19;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t20;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t21;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t22;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t23;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t24;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t25;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t26;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t27;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t28;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t29;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t30;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t31;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t32;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t33;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t34;
reg [2048-1:0] FSM_dct_8x8_stage_2_0_t35;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t36;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t37;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t38;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t39;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t40;
reg [2048-1:0] FSM_dct_8x8_stage_2_0_t41;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t42;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t43;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t44;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t45;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t46;
reg [2048-1:0] FSM_dct_8x8_stage_2_0_t47;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t48;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t49;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t50;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t51;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t52;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t53;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t54;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t55;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t56;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t57;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t58;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t59;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t60;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t61;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t62;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t63;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t64;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t65;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t66;
reg [2048-1:0] FSM_dct_8x8_stage_2_0_t67;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t68;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t69;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t70;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t71;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t72;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t73;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t74;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t75;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t76;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t77;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t78;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t79;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t80;
reg [2048-1:0] FSM_dct_8x8_stage_2_0_t81;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t82;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t83;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t84;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t85;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t86;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t87;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t88;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t89;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t90;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t91;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t92;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t93;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t94;
reg [2048-1:0] FSM_dct_8x8_stage_2_0_t95;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t96;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t97;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t98;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t99;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t100;
reg [2048-1:0] FSM_dct_8x8_stage_2_0_t101;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t102;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t103;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t104;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t105;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t106;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t107;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t108;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t109;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t110;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t111;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t112;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t113;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t114;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t115;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t116;
reg [2048-1:0] FSM_dct_8x8_stage_2_0_t117;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t118;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t119;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t120;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t121;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t122;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t123;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t124;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t125;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t126;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t127;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t128;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t129;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t130;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t131;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t132;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t133;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t134;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t135;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t136;
reg [2048-1:0] FSM_dct_8x8_stage_2_0_t137;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t138;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t139;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t140;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t141;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t142;
reg [2048-1:0] FSM_dct_8x8_stage_2_0_t143;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t144;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t145;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t146;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t147;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t148;
reg [2048-1:0] FSM_dct_8x8_stage_2_0_t149;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t150;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t151;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t152;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t153;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t154;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t155;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t156;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t157;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t158;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t159;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t160;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t161;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t162;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t163;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t164;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t165;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t166;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t167;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t168;
reg [2048-1:0] FSM_dct_8x8_stage_2_0_t169;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t170;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t171;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t172;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t173;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t174;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t175;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t176;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t177;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t178;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t179;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t180;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t181;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t182;
reg [2048-1:0] FSM_dct_8x8_stage_2_0_t183;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t184;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t185;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t186;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t187;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t188;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t189;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t190;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t191;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t192;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t193;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t194;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t195;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t196;
reg [2048-1:0] FSM_dct_8x8_stage_2_0_t197;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t198;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t199;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t200;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t201;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t202;
reg [2048-1:0] FSM_dct_8x8_stage_2_0_t203;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t204;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t205;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t206;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t207;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t208;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t209;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t210;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t211;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t212;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t213;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t214;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t215;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t216;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t217;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t218;
reg [2048-1:0] FSM_dct_8x8_stage_2_0_t219;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t220;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t221;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t222;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t223;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t224;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t225;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t226;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t227;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t228;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t229;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t230;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t231;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t232;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t233;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t234;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t235;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t236;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t237;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t238;
reg [2048-1:0] FSM_dct_8x8_stage_2_0_t239;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t240;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t241;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t242;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t243;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t244;
reg [2048-1:0] FSM_dct_8x8_stage_2_0_t245;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t246;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t247;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t248;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t249;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t250;
reg [2048-1:0] FSM_dct_8x8_stage_2_0_t251;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t252;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t253;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t254;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t255;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t256;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t257;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t258;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t259;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t260;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t261;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t262;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t263;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t264;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t265;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t266;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t267;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t268;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t269;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t270;
reg [2048-1:0] FSM_dct_8x8_stage_2_0_t271;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t272;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t273;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t274;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t275;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t276;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t277;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t278;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t279;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t280;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t281;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t282;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t283;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t284;
reg [2048-1:0] FSM_dct_8x8_stage_2_0_t285;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t286;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t287;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t288;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t289;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t290;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t291;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t292;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t293;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t294;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t295;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t296;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t297;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t298;
reg [2048-1:0] FSM_dct_8x8_stage_2_0_t299;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t300;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t301;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t302;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t303;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t304;
reg [2048-1:0] FSM_dct_8x8_stage_2_0_t305;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t306;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t307;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t308;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t309;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t310;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t311;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t312;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t313;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t314;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t315;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t316;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t317;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t318;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t319;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t320;
reg [2048-1:0] FSM_dct_8x8_stage_2_0_t321;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t322;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t323;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t324;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t325;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t326;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t327;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t328;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t329;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t330;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t331;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t332;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t333;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t334;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t335;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t336;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t337;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t338;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t339;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t340;
reg [2048-1:0] FSM_dct_8x8_stage_2_0_t341;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t342;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t343;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t344;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t345;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t346;
reg [2048-1:0] FSM_dct_8x8_stage_2_0_t347;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t348;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t349;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t350;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t351;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t352;
reg [2048-1:0] FSM_dct_8x8_stage_2_0_t353;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t354;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t355;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t356;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t357;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t358;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t359;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t360;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t361;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t362;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t363;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t364;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t365;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t366;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t367;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t368;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t369;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t370;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t371;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t372;
reg [2048-1:0] FSM_dct_8x8_stage_2_0_t373;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t374;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t375;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t376;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t377;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t378;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t379;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t380;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t381;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t382;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t383;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t384;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t385;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t386;
reg [2048-1:0] FSM_dct_8x8_stage_2_0_t387;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t388;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t389;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t390;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t391;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t392;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t393;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t394;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t395;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t396;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t397;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t398;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t399;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t400;
reg [2048-1:0] FSM_dct_8x8_stage_2_0_t401;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t402;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t403;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t404;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t405;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t406;
reg [2048-1:0] FSM_dct_8x8_stage_2_0_t407;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t408;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t409;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t410;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t411;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t412;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t413;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t414;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t415;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t416;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t417;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t418;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t419;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t420;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t421;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t422;
reg [2048-1:0] FSM_dct_8x8_stage_2_0_t423;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t424;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t425;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t426;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t427;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t428;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t429;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t430;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t431;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t432;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t433;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t434;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t435;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t436;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t437;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t438;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t439;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t440;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t441;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t442;
reg [2048-1:0] FSM_dct_8x8_stage_2_0_t443;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t444;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t445;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t446;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t447;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t448;
reg [2048-1:0] FSM_dct_8x8_stage_2_0_t449;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t450;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t451;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t452;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t453;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t454;
reg [2048-1:0] FSM_dct_8x8_stage_2_0_t455;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t456;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t457;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t458;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t459;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t460;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t461;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t462;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t463;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t464;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t465;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t466;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t467;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t468;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t469;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t470;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t471;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t472;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t473;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t474;
reg [2048-1:0] FSM_dct_8x8_stage_2_0_t475;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t476;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t477;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t478;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t479;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t480;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t481;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t482;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t483;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t484;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t485;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t486;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t487;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t488;
reg [2048-1:0] FSM_dct_8x8_stage_2_0_t489;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t490;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t491;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t492;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t493;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t494;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t495;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t496;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t497;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t498;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t499;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t500;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t501;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t502;
reg [2048-1:0] FSM_dct_8x8_stage_2_0_t503;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t504;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t505;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t506;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t507;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t508;
reg [2048-1:0] FSM_dct_8x8_stage_2_0_t509;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t510;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t511;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t512;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t513;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t514;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t515;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t516;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t517;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t518;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t519;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t520;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t521;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t522;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t523;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t524;
reg [2048-1:0] FSM_dct_8x8_stage_2_0_t525;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t526;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t527;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t528;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t529;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t530;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t531;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t532;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t533;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t534;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t535;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t536;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t537;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t538;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t539;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t540;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t541;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t542;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t543;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t544;
reg [2048-1:0] FSM_dct_8x8_stage_2_0_t545;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t546;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t547;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t548;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t549;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t550;
reg [2048-1:0] FSM_dct_8x8_stage_2_0_t551;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t552;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t553;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t554;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t555;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t556;
reg [2048-1:0] FSM_dct_8x8_stage_2_0_t557;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t558;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t559;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t560;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t561;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t562;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t563;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t564;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t565;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t566;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t567;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t568;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t569;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t570;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t571;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t572;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t573;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t574;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t575;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t576;
reg [2048-1:0] FSM_dct_8x8_stage_2_0_t577;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t578;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t579;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t580;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t581;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t582;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t583;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t584;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t585;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t586;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t587;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t588;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t589;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t590;
reg [2048-1:0] FSM_dct_8x8_stage_2_0_t591;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t592;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t593;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t594;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t595;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t596;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t597;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t598;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t599;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t600;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t601;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t602;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t603;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t604;
reg [2048-1:0] FSM_dct_8x8_stage_2_0_t605;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t606;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t607;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t608;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t609;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t610;
reg [2048-1:0] FSM_dct_8x8_stage_2_0_t611;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t612;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t613;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t614;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t615;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t616;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t617;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t618;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t619;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t620;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t621;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t622;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t623;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t624;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t625;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t626;
reg [2048-1:0] FSM_dct_8x8_stage_2_0_t627;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t628;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t629;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t630;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t631;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t632;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t633;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t634;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t635;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t636;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t637;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t638;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t639;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t640;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t641;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t642;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t643;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t644;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t645;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t646;
reg [2048-1:0] FSM_dct_8x8_stage_2_0_t647;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t648;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t649;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t650;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t651;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t652;
reg [2048-1:0] FSM_dct_8x8_stage_2_0_t653;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t654;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t655;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t656;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t657;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t658;
reg [2048-1:0] FSM_dct_8x8_stage_2_0_t659;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t660;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t661;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t662;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t663;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t664;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t665;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t666;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t667;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t668;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t669;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t670;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t671;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t672;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t673;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t674;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t675;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t676;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t677;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t678;
reg [2048-1:0] FSM_dct_8x8_stage_2_0_t679;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t680;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t681;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t682;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t683;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t684;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t685;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t686;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t687;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t688;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t689;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t690;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t691;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t692;
reg [2048-1:0] FSM_dct_8x8_stage_2_0_t693;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t694;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t695;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t696;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t697;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t698;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t699;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t700;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t701;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t702;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t703;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t704;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t705;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t706;
reg [2048-1:0] FSM_dct_8x8_stage_2_0_t707;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t708;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t709;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t710;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t711;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t712;
reg [2048-1:0] FSM_dct_8x8_stage_2_0_t713;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t714;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t715;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t716;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t717;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t718;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t719;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t720;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t721;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t722;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t723;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t724;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t725;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t726;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t727;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t728;
reg [2048-1:0] FSM_dct_8x8_stage_2_0_t729;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t730;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t731;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t732;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t733;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t734;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t735;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t736;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t737;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t738;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t739;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t740;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t741;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t742;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t743;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t744;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t745;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t746;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t747;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t748;
reg [2048-1:0] FSM_dct_8x8_stage_2_0_t749;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t750;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t751;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t752;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t753;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t754;
reg [2048-1:0] FSM_dct_8x8_stage_2_0_t755;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t756;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t757;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t758;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t759;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t760;
reg [2048-1:0] FSM_dct_8x8_stage_2_0_t761;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t762;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t763;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t764;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t765;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t766;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t767;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t768;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t769;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t770;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t771;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t772;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t773;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t774;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t775;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t776;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t777;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t778;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t779;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t780;
reg [2048-1:0] FSM_dct_8x8_stage_2_0_t781;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t782;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t783;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t784;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t785;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t786;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t787;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t788;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t789;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t790;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t791;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t792;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t793;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t794;
reg [2048-1:0] FSM_dct_8x8_stage_2_0_t795;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t796;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t797;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t798;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t799;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t800;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t801;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t802;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t803;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t804;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t805;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t806;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t807;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t808;
reg [2048-1:0] FSM_dct_8x8_stage_2_0_t809;
reg [64-1:0] FSM_dct_8x8_stage_2_0_t810;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t811;
reg [33-1:0] FSM_dct_8x8_stage_2_0_t812;
reg [32-1:0] FSM_dct_8x8_stage_2_0_t813;
reg [6-1:0] FSM_dct_8x8_stage_2_0_t814;
reg [2048-1:0] FSM_dct_8x8_stage_2_0_t815;

/*
    Wiring by dct_8x8_stage_2
*/
assign i_ready = FSM_dct_8x8_stage_2_0_in_ready;
assign o_data_out = FSM_dct_8x8_stage_2_0_t815;
assign o_valid = FSM_dct_8x8_stage_2_0_out_valid;
/* End wiring by dct_8x8_stage_2 */

assign FSM_dct_8x8_stage_2_0_out_valid = 1'b1;

initial begin
    FSM_dct_8x8_stage_2_0_t0 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_2_0_t1 = FSM_dct_8x8_stage_2_0_t0[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t2 = FSM_dct_8x8_stage_2_0_t1[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t3 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_2_0_t4 = FSM_dct_8x8_stage_2_0_t3[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t5 = FSM_dct_8x8_stage_2_0_t4[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t6 = i_data_in[FSM_dct_8x8_stage_2_0_t5 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t7 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_2_0_t8 = FSM_dct_8x8_stage_2_0_t7[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t9 = FSM_dct_8x8_stage_2_0_t8 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_2_0_t10 = FSM_dct_8x8_stage_2_0_t9[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t11 = FSM_dct_8x8_stage_2_0_t10[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t12 = i_data_in[FSM_dct_8x8_stage_2_0_t11 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t13 = FSM_dct_8x8_stage_2_0_t6 + FSM_dct_8x8_stage_2_0_t12;
    FSM_dct_8x8_stage_2_0_t14 = FSM_dct_8x8_stage_2_0_t13[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t15 = 2048'b0;
    FSM_dct_8x8_stage_2_0_t15[FSM_dct_8x8_stage_2_0_t2 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t14;
    FSM_dct_8x8_stage_2_0_t16 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_2_0_t17 = FSM_dct_8x8_stage_2_0_t16[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t18 = FSM_dct_8x8_stage_2_0_t17 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_2_0_t19 = FSM_dct_8x8_stage_2_0_t18[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t20 = FSM_dct_8x8_stage_2_0_t19[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t21 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_2_0_t22 = FSM_dct_8x8_stage_2_0_t21[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t23 = FSM_dct_8x8_stage_2_0_t22 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_2_0_t24 = FSM_dct_8x8_stage_2_0_t23[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t25 = FSM_dct_8x8_stage_2_0_t24[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t26 = i_data_in[FSM_dct_8x8_stage_2_0_t25 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t27 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_2_0_t28 = FSM_dct_8x8_stage_2_0_t27[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t29 = FSM_dct_8x8_stage_2_0_t28 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_2_0_t30 = FSM_dct_8x8_stage_2_0_t29[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t31 = FSM_dct_8x8_stage_2_0_t30[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t32 = i_data_in[FSM_dct_8x8_stage_2_0_t31 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t33 = FSM_dct_8x8_stage_2_0_t26 + FSM_dct_8x8_stage_2_0_t32;
    FSM_dct_8x8_stage_2_0_t34 = FSM_dct_8x8_stage_2_0_t33[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t35 = FSM_dct_8x8_stage_2_0_t15;
    FSM_dct_8x8_stage_2_0_t35[FSM_dct_8x8_stage_2_0_t20 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t34;
    FSM_dct_8x8_stage_2_0_t36 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_2_0_t37 = FSM_dct_8x8_stage_2_0_t36[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t38 = FSM_dct_8x8_stage_2_0_t37 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_2_0_t39 = FSM_dct_8x8_stage_2_0_t38[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t40 = FSM_dct_8x8_stage_2_0_t39[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t41 = FSM_dct_8x8_stage_2_0_t35;
    FSM_dct_8x8_stage_2_0_t41[FSM_dct_8x8_stage_2_0_t40 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t26 - FSM_dct_8x8_stage_2_0_t32;
    FSM_dct_8x8_stage_2_0_t42 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_2_0_t43 = FSM_dct_8x8_stage_2_0_t42[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t44 = FSM_dct_8x8_stage_2_0_t43 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_2_0_t45 = FSM_dct_8x8_stage_2_0_t44[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t46 = FSM_dct_8x8_stage_2_0_t45[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t47 = FSM_dct_8x8_stage_2_0_t41;
    FSM_dct_8x8_stage_2_0_t47[FSM_dct_8x8_stage_2_0_t46 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t6 - FSM_dct_8x8_stage_2_0_t12;
    FSM_dct_8x8_stage_2_0_t48 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_2_0_t49 = FSM_dct_8x8_stage_2_0_t48[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t50 = FSM_dct_8x8_stage_2_0_t49 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_2_0_t51 = FSM_dct_8x8_stage_2_0_t50[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t52 = FSM_dct_8x8_stage_2_0_t51[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t53 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_2_0_t54 = FSM_dct_8x8_stage_2_0_t53[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t55 = FSM_dct_8x8_stage_2_0_t54 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_2_0_t56 = FSM_dct_8x8_stage_2_0_t55[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t57 = FSM_dct_8x8_stage_2_0_t56[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t58 = i_data_in[FSM_dct_8x8_stage_2_0_t57 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t59 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_2_0_t60 = FSM_dct_8x8_stage_2_0_t59[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t61 = FSM_dct_8x8_stage_2_0_t60 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_2_0_t62 = FSM_dct_8x8_stage_2_0_t61[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t63 = FSM_dct_8x8_stage_2_0_t62[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t64 = i_data_in[FSM_dct_8x8_stage_2_0_t63 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t65 = FSM_dct_8x8_stage_2_0_t58 + FSM_dct_8x8_stage_2_0_t64;
    FSM_dct_8x8_stage_2_0_t66 = FSM_dct_8x8_stage_2_0_t65[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t67 = FSM_dct_8x8_stage_2_0_t47;
    FSM_dct_8x8_stage_2_0_t67[FSM_dct_8x8_stage_2_0_t52 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t66;
    FSM_dct_8x8_stage_2_0_t68 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_2_0_t69 = FSM_dct_8x8_stage_2_0_t68[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t70 = FSM_dct_8x8_stage_2_0_t69 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_2_0_t71 = FSM_dct_8x8_stage_2_0_t70[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t72 = FSM_dct_8x8_stage_2_0_t71[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t73 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_2_0_t74 = FSM_dct_8x8_stage_2_0_t73[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t75 = FSM_dct_8x8_stage_2_0_t74 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_2_0_t76 = FSM_dct_8x8_stage_2_0_t75[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t77 = FSM_dct_8x8_stage_2_0_t76[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t78 = i_data_in[FSM_dct_8x8_stage_2_0_t77 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t79 = FSM_dct_8x8_stage_2_0_t64 + FSM_dct_8x8_stage_2_0_t78;
    FSM_dct_8x8_stage_2_0_t80 = FSM_dct_8x8_stage_2_0_t79[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t81 = FSM_dct_8x8_stage_2_0_t67;
    FSM_dct_8x8_stage_2_0_t81[FSM_dct_8x8_stage_2_0_t72 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t80;
    FSM_dct_8x8_stage_2_0_t82 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_2_0_t83 = FSM_dct_8x8_stage_2_0_t82[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t84 = FSM_dct_8x8_stage_2_0_t83 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_2_0_t85 = FSM_dct_8x8_stage_2_0_t84[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t86 = FSM_dct_8x8_stage_2_0_t85[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t87 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_2_0_t88 = FSM_dct_8x8_stage_2_0_t87[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t89 = FSM_dct_8x8_stage_2_0_t88 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_2_0_t90 = FSM_dct_8x8_stage_2_0_t89[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t91 = FSM_dct_8x8_stage_2_0_t90[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t92 = i_data_in[FSM_dct_8x8_stage_2_0_t91 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t93 = FSM_dct_8x8_stage_2_0_t78 + FSM_dct_8x8_stage_2_0_t92;
    FSM_dct_8x8_stage_2_0_t94 = FSM_dct_8x8_stage_2_0_t93[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t95 = FSM_dct_8x8_stage_2_0_t81;
    FSM_dct_8x8_stage_2_0_t95[FSM_dct_8x8_stage_2_0_t86 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t94;
    FSM_dct_8x8_stage_2_0_t96 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_2_0_t97 = FSM_dct_8x8_stage_2_0_t96[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t98 = FSM_dct_8x8_stage_2_0_t97 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_2_0_t99 = FSM_dct_8x8_stage_2_0_t98[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t100 = FSM_dct_8x8_stage_2_0_t99[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t101 = FSM_dct_8x8_stage_2_0_t95;
    FSM_dct_8x8_stage_2_0_t101[FSM_dct_8x8_stage_2_0_t100 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t92;
    FSM_dct_8x8_stage_2_0_t102 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_2_0_t103 = FSM_dct_8x8_stage_2_0_t102[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t104 = FSM_dct_8x8_stage_2_0_t103[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t105 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_2_0_t106 = FSM_dct_8x8_stage_2_0_t105[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t107 = FSM_dct_8x8_stage_2_0_t106[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t108 = i_data_in[FSM_dct_8x8_stage_2_0_t107 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t109 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_2_0_t110 = FSM_dct_8x8_stage_2_0_t109[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t111 = FSM_dct_8x8_stage_2_0_t110 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_2_0_t112 = FSM_dct_8x8_stage_2_0_t111[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t113 = FSM_dct_8x8_stage_2_0_t112[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t114 = i_data_in[FSM_dct_8x8_stage_2_0_t113 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t115 = FSM_dct_8x8_stage_2_0_t108 + FSM_dct_8x8_stage_2_0_t114;
    FSM_dct_8x8_stage_2_0_t116 = FSM_dct_8x8_stage_2_0_t115[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t117 = FSM_dct_8x8_stage_2_0_t101;
    FSM_dct_8x8_stage_2_0_t117[FSM_dct_8x8_stage_2_0_t104 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t116;
    FSM_dct_8x8_stage_2_0_t118 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_2_0_t119 = FSM_dct_8x8_stage_2_0_t118[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t120 = FSM_dct_8x8_stage_2_0_t119 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_2_0_t121 = FSM_dct_8x8_stage_2_0_t120[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t122 = FSM_dct_8x8_stage_2_0_t121[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t123 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_2_0_t124 = FSM_dct_8x8_stage_2_0_t123[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t125 = FSM_dct_8x8_stage_2_0_t124 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_2_0_t126 = FSM_dct_8x8_stage_2_0_t125[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t127 = FSM_dct_8x8_stage_2_0_t126[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t128 = i_data_in[FSM_dct_8x8_stage_2_0_t127 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t129 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_2_0_t130 = FSM_dct_8x8_stage_2_0_t129[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t131 = FSM_dct_8x8_stage_2_0_t130 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_2_0_t132 = FSM_dct_8x8_stage_2_0_t131[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t133 = FSM_dct_8x8_stage_2_0_t132[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t134 = i_data_in[FSM_dct_8x8_stage_2_0_t133 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t135 = FSM_dct_8x8_stage_2_0_t128 + FSM_dct_8x8_stage_2_0_t134;
    FSM_dct_8x8_stage_2_0_t136 = FSM_dct_8x8_stage_2_0_t135[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t137 = FSM_dct_8x8_stage_2_0_t117;
    FSM_dct_8x8_stage_2_0_t137[FSM_dct_8x8_stage_2_0_t122 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t136;
    FSM_dct_8x8_stage_2_0_t138 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_2_0_t139 = FSM_dct_8x8_stage_2_0_t138[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t140 = FSM_dct_8x8_stage_2_0_t139 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_2_0_t141 = FSM_dct_8x8_stage_2_0_t140[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t142 = FSM_dct_8x8_stage_2_0_t141[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t143 = FSM_dct_8x8_stage_2_0_t137;
    FSM_dct_8x8_stage_2_0_t143[FSM_dct_8x8_stage_2_0_t142 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t128 - FSM_dct_8x8_stage_2_0_t134;
    FSM_dct_8x8_stage_2_0_t144 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_2_0_t145 = FSM_dct_8x8_stage_2_0_t144[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t146 = FSM_dct_8x8_stage_2_0_t145 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_2_0_t147 = FSM_dct_8x8_stage_2_0_t146[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t148 = FSM_dct_8x8_stage_2_0_t147[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t149 = FSM_dct_8x8_stage_2_0_t143;
    FSM_dct_8x8_stage_2_0_t149[FSM_dct_8x8_stage_2_0_t148 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t108 - FSM_dct_8x8_stage_2_0_t114;
    FSM_dct_8x8_stage_2_0_t150 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_2_0_t151 = FSM_dct_8x8_stage_2_0_t150[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t152 = FSM_dct_8x8_stage_2_0_t151 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_2_0_t153 = FSM_dct_8x8_stage_2_0_t152[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t154 = FSM_dct_8x8_stage_2_0_t153[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t155 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_2_0_t156 = FSM_dct_8x8_stage_2_0_t155[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t157 = FSM_dct_8x8_stage_2_0_t156 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_2_0_t158 = FSM_dct_8x8_stage_2_0_t157[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t159 = FSM_dct_8x8_stage_2_0_t158[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t160 = i_data_in[FSM_dct_8x8_stage_2_0_t159 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t161 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_2_0_t162 = FSM_dct_8x8_stage_2_0_t161[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t163 = FSM_dct_8x8_stage_2_0_t162 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_2_0_t164 = FSM_dct_8x8_stage_2_0_t163[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t165 = FSM_dct_8x8_stage_2_0_t164[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t166 = i_data_in[FSM_dct_8x8_stage_2_0_t165 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t167 = FSM_dct_8x8_stage_2_0_t160 + FSM_dct_8x8_stage_2_0_t166;
    FSM_dct_8x8_stage_2_0_t168 = FSM_dct_8x8_stage_2_0_t167[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t169 = FSM_dct_8x8_stage_2_0_t149;
    FSM_dct_8x8_stage_2_0_t169[FSM_dct_8x8_stage_2_0_t154 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t168;
    FSM_dct_8x8_stage_2_0_t170 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_2_0_t171 = FSM_dct_8x8_stage_2_0_t170[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t172 = FSM_dct_8x8_stage_2_0_t171 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_2_0_t173 = FSM_dct_8x8_stage_2_0_t172[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t174 = FSM_dct_8x8_stage_2_0_t173[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t175 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_2_0_t176 = FSM_dct_8x8_stage_2_0_t175[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t177 = FSM_dct_8x8_stage_2_0_t176 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_2_0_t178 = FSM_dct_8x8_stage_2_0_t177[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t179 = FSM_dct_8x8_stage_2_0_t178[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t180 = i_data_in[FSM_dct_8x8_stage_2_0_t179 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t181 = FSM_dct_8x8_stage_2_0_t166 + FSM_dct_8x8_stage_2_0_t180;
    FSM_dct_8x8_stage_2_0_t182 = FSM_dct_8x8_stage_2_0_t181[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t183 = FSM_dct_8x8_stage_2_0_t169;
    FSM_dct_8x8_stage_2_0_t183[FSM_dct_8x8_stage_2_0_t174 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t182;
    FSM_dct_8x8_stage_2_0_t184 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_2_0_t185 = FSM_dct_8x8_stage_2_0_t184[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t186 = FSM_dct_8x8_stage_2_0_t185 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_2_0_t187 = FSM_dct_8x8_stage_2_0_t186[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t188 = FSM_dct_8x8_stage_2_0_t187[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t189 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_2_0_t190 = FSM_dct_8x8_stage_2_0_t189[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t191 = FSM_dct_8x8_stage_2_0_t190 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_2_0_t192 = FSM_dct_8x8_stage_2_0_t191[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t193 = FSM_dct_8x8_stage_2_0_t192[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t194 = i_data_in[FSM_dct_8x8_stage_2_0_t193 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t195 = FSM_dct_8x8_stage_2_0_t180 + FSM_dct_8x8_stage_2_0_t194;
    FSM_dct_8x8_stage_2_0_t196 = FSM_dct_8x8_stage_2_0_t195[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t197 = FSM_dct_8x8_stage_2_0_t183;
    FSM_dct_8x8_stage_2_0_t197[FSM_dct_8x8_stage_2_0_t188 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t196;
    FSM_dct_8x8_stage_2_0_t198 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_2_0_t199 = FSM_dct_8x8_stage_2_0_t198[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t200 = FSM_dct_8x8_stage_2_0_t199 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_2_0_t201 = FSM_dct_8x8_stage_2_0_t200[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t202 = FSM_dct_8x8_stage_2_0_t201[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t203 = FSM_dct_8x8_stage_2_0_t197;
    FSM_dct_8x8_stage_2_0_t203[FSM_dct_8x8_stage_2_0_t202 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t194;
    FSM_dct_8x8_stage_2_0_t204 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_2_0_t205 = FSM_dct_8x8_stage_2_0_t204[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t206 = FSM_dct_8x8_stage_2_0_t205[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t207 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_2_0_t208 = FSM_dct_8x8_stage_2_0_t207[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t209 = FSM_dct_8x8_stage_2_0_t208[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t210 = i_data_in[FSM_dct_8x8_stage_2_0_t209 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t211 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_2_0_t212 = FSM_dct_8x8_stage_2_0_t211[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t213 = FSM_dct_8x8_stage_2_0_t212 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_2_0_t214 = FSM_dct_8x8_stage_2_0_t213[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t215 = FSM_dct_8x8_stage_2_0_t214[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t216 = i_data_in[FSM_dct_8x8_stage_2_0_t215 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t217 = FSM_dct_8x8_stage_2_0_t210 + FSM_dct_8x8_stage_2_0_t216;
    FSM_dct_8x8_stage_2_0_t218 = FSM_dct_8x8_stage_2_0_t217[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t219 = FSM_dct_8x8_stage_2_0_t203;
    FSM_dct_8x8_stage_2_0_t219[FSM_dct_8x8_stage_2_0_t206 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t218;
    FSM_dct_8x8_stage_2_0_t220 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_2_0_t221 = FSM_dct_8x8_stage_2_0_t220[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t222 = FSM_dct_8x8_stage_2_0_t221 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_2_0_t223 = FSM_dct_8x8_stage_2_0_t222[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t224 = FSM_dct_8x8_stage_2_0_t223[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t225 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_2_0_t226 = FSM_dct_8x8_stage_2_0_t225[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t227 = FSM_dct_8x8_stage_2_0_t226 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_2_0_t228 = FSM_dct_8x8_stage_2_0_t227[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t229 = FSM_dct_8x8_stage_2_0_t228[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t230 = i_data_in[FSM_dct_8x8_stage_2_0_t229 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t231 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_2_0_t232 = FSM_dct_8x8_stage_2_0_t231[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t233 = FSM_dct_8x8_stage_2_0_t232 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_2_0_t234 = FSM_dct_8x8_stage_2_0_t233[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t235 = FSM_dct_8x8_stage_2_0_t234[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t236 = i_data_in[FSM_dct_8x8_stage_2_0_t235 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t237 = FSM_dct_8x8_stage_2_0_t230 + FSM_dct_8x8_stage_2_0_t236;
    FSM_dct_8x8_stage_2_0_t238 = FSM_dct_8x8_stage_2_0_t237[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t239 = FSM_dct_8x8_stage_2_0_t219;
    FSM_dct_8x8_stage_2_0_t239[FSM_dct_8x8_stage_2_0_t224 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t238;
    FSM_dct_8x8_stage_2_0_t240 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_2_0_t241 = FSM_dct_8x8_stage_2_0_t240[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t242 = FSM_dct_8x8_stage_2_0_t241 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_2_0_t243 = FSM_dct_8x8_stage_2_0_t242[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t244 = FSM_dct_8x8_stage_2_0_t243[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t245 = FSM_dct_8x8_stage_2_0_t239;
    FSM_dct_8x8_stage_2_0_t245[FSM_dct_8x8_stage_2_0_t244 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t230 - FSM_dct_8x8_stage_2_0_t236;
    FSM_dct_8x8_stage_2_0_t246 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_2_0_t247 = FSM_dct_8x8_stage_2_0_t246[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t248 = FSM_dct_8x8_stage_2_0_t247 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_2_0_t249 = FSM_dct_8x8_stage_2_0_t248[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t250 = FSM_dct_8x8_stage_2_0_t249[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t251 = FSM_dct_8x8_stage_2_0_t245;
    FSM_dct_8x8_stage_2_0_t251[FSM_dct_8x8_stage_2_0_t250 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t210 - FSM_dct_8x8_stage_2_0_t216;
    FSM_dct_8x8_stage_2_0_t252 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_2_0_t253 = FSM_dct_8x8_stage_2_0_t252[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t254 = FSM_dct_8x8_stage_2_0_t253 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_2_0_t255 = FSM_dct_8x8_stage_2_0_t254[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t256 = FSM_dct_8x8_stage_2_0_t255[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t257 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_2_0_t258 = FSM_dct_8x8_stage_2_0_t257[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t259 = FSM_dct_8x8_stage_2_0_t258 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_2_0_t260 = FSM_dct_8x8_stage_2_0_t259[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t261 = FSM_dct_8x8_stage_2_0_t260[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t262 = i_data_in[FSM_dct_8x8_stage_2_0_t261 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t263 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_2_0_t264 = FSM_dct_8x8_stage_2_0_t263[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t265 = FSM_dct_8x8_stage_2_0_t264 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_2_0_t266 = FSM_dct_8x8_stage_2_0_t265[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t267 = FSM_dct_8x8_stage_2_0_t266[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t268 = i_data_in[FSM_dct_8x8_stage_2_0_t267 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t269 = FSM_dct_8x8_stage_2_0_t262 + FSM_dct_8x8_stage_2_0_t268;
    FSM_dct_8x8_stage_2_0_t270 = FSM_dct_8x8_stage_2_0_t269[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t271 = FSM_dct_8x8_stage_2_0_t251;
    FSM_dct_8x8_stage_2_0_t271[FSM_dct_8x8_stage_2_0_t256 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t270;
    FSM_dct_8x8_stage_2_0_t272 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_2_0_t273 = FSM_dct_8x8_stage_2_0_t272[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t274 = FSM_dct_8x8_stage_2_0_t273 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_2_0_t275 = FSM_dct_8x8_stage_2_0_t274[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t276 = FSM_dct_8x8_stage_2_0_t275[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t277 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_2_0_t278 = FSM_dct_8x8_stage_2_0_t277[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t279 = FSM_dct_8x8_stage_2_0_t278 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_2_0_t280 = FSM_dct_8x8_stage_2_0_t279[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t281 = FSM_dct_8x8_stage_2_0_t280[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t282 = i_data_in[FSM_dct_8x8_stage_2_0_t281 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t283 = FSM_dct_8x8_stage_2_0_t268 + FSM_dct_8x8_stage_2_0_t282;
    FSM_dct_8x8_stage_2_0_t284 = FSM_dct_8x8_stage_2_0_t283[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t285 = FSM_dct_8x8_stage_2_0_t271;
    FSM_dct_8x8_stage_2_0_t285[FSM_dct_8x8_stage_2_0_t276 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t284;
    FSM_dct_8x8_stage_2_0_t286 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_2_0_t287 = FSM_dct_8x8_stage_2_0_t286[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t288 = FSM_dct_8x8_stage_2_0_t287 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_2_0_t289 = FSM_dct_8x8_stage_2_0_t288[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t290 = FSM_dct_8x8_stage_2_0_t289[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t291 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_2_0_t292 = FSM_dct_8x8_stage_2_0_t291[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t293 = FSM_dct_8x8_stage_2_0_t292 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_2_0_t294 = FSM_dct_8x8_stage_2_0_t293[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t295 = FSM_dct_8x8_stage_2_0_t294[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t296 = i_data_in[FSM_dct_8x8_stage_2_0_t295 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t297 = FSM_dct_8x8_stage_2_0_t282 + FSM_dct_8x8_stage_2_0_t296;
    FSM_dct_8x8_stage_2_0_t298 = FSM_dct_8x8_stage_2_0_t297[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t299 = FSM_dct_8x8_stage_2_0_t285;
    FSM_dct_8x8_stage_2_0_t299[FSM_dct_8x8_stage_2_0_t290 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t298;
    FSM_dct_8x8_stage_2_0_t300 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_2_0_t301 = FSM_dct_8x8_stage_2_0_t300[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t302 = FSM_dct_8x8_stage_2_0_t301 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_2_0_t303 = FSM_dct_8x8_stage_2_0_t302[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t304 = FSM_dct_8x8_stage_2_0_t303[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t305 = FSM_dct_8x8_stage_2_0_t299;
    FSM_dct_8x8_stage_2_0_t305[FSM_dct_8x8_stage_2_0_t304 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t296;
    FSM_dct_8x8_stage_2_0_t306 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_2_0_t307 = FSM_dct_8x8_stage_2_0_t306[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t308 = FSM_dct_8x8_stage_2_0_t307[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t309 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_2_0_t310 = FSM_dct_8x8_stage_2_0_t309[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t311 = FSM_dct_8x8_stage_2_0_t310[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t312 = i_data_in[FSM_dct_8x8_stage_2_0_t311 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t313 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_2_0_t314 = FSM_dct_8x8_stage_2_0_t313[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t315 = FSM_dct_8x8_stage_2_0_t314 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_2_0_t316 = FSM_dct_8x8_stage_2_0_t315[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t317 = FSM_dct_8x8_stage_2_0_t316[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t318 = i_data_in[FSM_dct_8x8_stage_2_0_t317 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t319 = FSM_dct_8x8_stage_2_0_t312 + FSM_dct_8x8_stage_2_0_t318;
    FSM_dct_8x8_stage_2_0_t320 = FSM_dct_8x8_stage_2_0_t319[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t321 = FSM_dct_8x8_stage_2_0_t305;
    FSM_dct_8x8_stage_2_0_t321[FSM_dct_8x8_stage_2_0_t308 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t320;
    FSM_dct_8x8_stage_2_0_t322 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_2_0_t323 = FSM_dct_8x8_stage_2_0_t322[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t324 = FSM_dct_8x8_stage_2_0_t323 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_2_0_t325 = FSM_dct_8x8_stage_2_0_t324[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t326 = FSM_dct_8x8_stage_2_0_t325[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t327 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_2_0_t328 = FSM_dct_8x8_stage_2_0_t327[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t329 = FSM_dct_8x8_stage_2_0_t328 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_2_0_t330 = FSM_dct_8x8_stage_2_0_t329[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t331 = FSM_dct_8x8_stage_2_0_t330[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t332 = i_data_in[FSM_dct_8x8_stage_2_0_t331 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t333 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_2_0_t334 = FSM_dct_8x8_stage_2_0_t333[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t335 = FSM_dct_8x8_stage_2_0_t334 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_2_0_t336 = FSM_dct_8x8_stage_2_0_t335[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t337 = FSM_dct_8x8_stage_2_0_t336[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t338 = i_data_in[FSM_dct_8x8_stage_2_0_t337 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t339 = FSM_dct_8x8_stage_2_0_t332 + FSM_dct_8x8_stage_2_0_t338;
    FSM_dct_8x8_stage_2_0_t340 = FSM_dct_8x8_stage_2_0_t339[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t341 = FSM_dct_8x8_stage_2_0_t321;
    FSM_dct_8x8_stage_2_0_t341[FSM_dct_8x8_stage_2_0_t326 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t340;
    FSM_dct_8x8_stage_2_0_t342 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_2_0_t343 = FSM_dct_8x8_stage_2_0_t342[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t344 = FSM_dct_8x8_stage_2_0_t343 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_2_0_t345 = FSM_dct_8x8_stage_2_0_t344[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t346 = FSM_dct_8x8_stage_2_0_t345[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t347 = FSM_dct_8x8_stage_2_0_t341;
    FSM_dct_8x8_stage_2_0_t347[FSM_dct_8x8_stage_2_0_t346 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t332 - FSM_dct_8x8_stage_2_0_t338;
    FSM_dct_8x8_stage_2_0_t348 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_2_0_t349 = FSM_dct_8x8_stage_2_0_t348[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t350 = FSM_dct_8x8_stage_2_0_t349 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_2_0_t351 = FSM_dct_8x8_stage_2_0_t350[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t352 = FSM_dct_8x8_stage_2_0_t351[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t353 = FSM_dct_8x8_stage_2_0_t347;
    FSM_dct_8x8_stage_2_0_t353[FSM_dct_8x8_stage_2_0_t352 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t312 - FSM_dct_8x8_stage_2_0_t318;
    FSM_dct_8x8_stage_2_0_t354 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_2_0_t355 = FSM_dct_8x8_stage_2_0_t354[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t356 = FSM_dct_8x8_stage_2_0_t355 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_2_0_t357 = FSM_dct_8x8_stage_2_0_t356[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t358 = FSM_dct_8x8_stage_2_0_t357[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t359 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_2_0_t360 = FSM_dct_8x8_stage_2_0_t359[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t361 = FSM_dct_8x8_stage_2_0_t360 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_2_0_t362 = FSM_dct_8x8_stage_2_0_t361[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t363 = FSM_dct_8x8_stage_2_0_t362[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t364 = i_data_in[FSM_dct_8x8_stage_2_0_t363 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t365 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_2_0_t366 = FSM_dct_8x8_stage_2_0_t365[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t367 = FSM_dct_8x8_stage_2_0_t366 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_2_0_t368 = FSM_dct_8x8_stage_2_0_t367[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t369 = FSM_dct_8x8_stage_2_0_t368[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t370 = i_data_in[FSM_dct_8x8_stage_2_0_t369 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t371 = FSM_dct_8x8_stage_2_0_t364 + FSM_dct_8x8_stage_2_0_t370;
    FSM_dct_8x8_stage_2_0_t372 = FSM_dct_8x8_stage_2_0_t371[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t373 = FSM_dct_8x8_stage_2_0_t353;
    FSM_dct_8x8_stage_2_0_t373[FSM_dct_8x8_stage_2_0_t358 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t372;
    FSM_dct_8x8_stage_2_0_t374 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_2_0_t375 = FSM_dct_8x8_stage_2_0_t374[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t376 = FSM_dct_8x8_stage_2_0_t375 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_2_0_t377 = FSM_dct_8x8_stage_2_0_t376[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t378 = FSM_dct_8x8_stage_2_0_t377[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t379 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_2_0_t380 = FSM_dct_8x8_stage_2_0_t379[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t381 = FSM_dct_8x8_stage_2_0_t380 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_2_0_t382 = FSM_dct_8x8_stage_2_0_t381[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t383 = FSM_dct_8x8_stage_2_0_t382[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t384 = i_data_in[FSM_dct_8x8_stage_2_0_t383 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t385 = FSM_dct_8x8_stage_2_0_t370 + FSM_dct_8x8_stage_2_0_t384;
    FSM_dct_8x8_stage_2_0_t386 = FSM_dct_8x8_stage_2_0_t385[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t387 = FSM_dct_8x8_stage_2_0_t373;
    FSM_dct_8x8_stage_2_0_t387[FSM_dct_8x8_stage_2_0_t378 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t386;
    FSM_dct_8x8_stage_2_0_t388 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_2_0_t389 = FSM_dct_8x8_stage_2_0_t388[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t390 = FSM_dct_8x8_stage_2_0_t389 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_2_0_t391 = FSM_dct_8x8_stage_2_0_t390[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t392 = FSM_dct_8x8_stage_2_0_t391[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t393 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_2_0_t394 = FSM_dct_8x8_stage_2_0_t393[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t395 = FSM_dct_8x8_stage_2_0_t394 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_2_0_t396 = FSM_dct_8x8_stage_2_0_t395[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t397 = FSM_dct_8x8_stage_2_0_t396[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t398 = i_data_in[FSM_dct_8x8_stage_2_0_t397 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t399 = FSM_dct_8x8_stage_2_0_t384 + FSM_dct_8x8_stage_2_0_t398;
    FSM_dct_8x8_stage_2_0_t400 = FSM_dct_8x8_stage_2_0_t399[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t401 = FSM_dct_8x8_stage_2_0_t387;
    FSM_dct_8x8_stage_2_0_t401[FSM_dct_8x8_stage_2_0_t392 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t400;
    FSM_dct_8x8_stage_2_0_t402 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_2_0_t403 = FSM_dct_8x8_stage_2_0_t402[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t404 = FSM_dct_8x8_stage_2_0_t403 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_2_0_t405 = FSM_dct_8x8_stage_2_0_t404[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t406 = FSM_dct_8x8_stage_2_0_t405[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t407 = FSM_dct_8x8_stage_2_0_t401;
    FSM_dct_8x8_stage_2_0_t407[FSM_dct_8x8_stage_2_0_t406 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t398;
    FSM_dct_8x8_stage_2_0_t408 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_2_0_t409 = FSM_dct_8x8_stage_2_0_t408[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t410 = FSM_dct_8x8_stage_2_0_t409[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t411 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_2_0_t412 = FSM_dct_8x8_stage_2_0_t411[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t413 = FSM_dct_8x8_stage_2_0_t412[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t414 = i_data_in[FSM_dct_8x8_stage_2_0_t413 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t415 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_2_0_t416 = FSM_dct_8x8_stage_2_0_t415[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t417 = FSM_dct_8x8_stage_2_0_t416 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_2_0_t418 = FSM_dct_8x8_stage_2_0_t417[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t419 = FSM_dct_8x8_stage_2_0_t418[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t420 = i_data_in[FSM_dct_8x8_stage_2_0_t419 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t421 = FSM_dct_8x8_stage_2_0_t414 + FSM_dct_8x8_stage_2_0_t420;
    FSM_dct_8x8_stage_2_0_t422 = FSM_dct_8x8_stage_2_0_t421[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t423 = FSM_dct_8x8_stage_2_0_t407;
    FSM_dct_8x8_stage_2_0_t423[FSM_dct_8x8_stage_2_0_t410 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t422;
    FSM_dct_8x8_stage_2_0_t424 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_2_0_t425 = FSM_dct_8x8_stage_2_0_t424[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t426 = FSM_dct_8x8_stage_2_0_t425 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_2_0_t427 = FSM_dct_8x8_stage_2_0_t426[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t428 = FSM_dct_8x8_stage_2_0_t427[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t429 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_2_0_t430 = FSM_dct_8x8_stage_2_0_t429[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t431 = FSM_dct_8x8_stage_2_0_t430 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_2_0_t432 = FSM_dct_8x8_stage_2_0_t431[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t433 = FSM_dct_8x8_stage_2_0_t432[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t434 = i_data_in[FSM_dct_8x8_stage_2_0_t433 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t435 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_2_0_t436 = FSM_dct_8x8_stage_2_0_t435[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t437 = FSM_dct_8x8_stage_2_0_t436 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_2_0_t438 = FSM_dct_8x8_stage_2_0_t437[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t439 = FSM_dct_8x8_stage_2_0_t438[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t440 = i_data_in[FSM_dct_8x8_stage_2_0_t439 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t441 = FSM_dct_8x8_stage_2_0_t434 + FSM_dct_8x8_stage_2_0_t440;
    FSM_dct_8x8_stage_2_0_t442 = FSM_dct_8x8_stage_2_0_t441[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t443 = FSM_dct_8x8_stage_2_0_t423;
    FSM_dct_8x8_stage_2_0_t443[FSM_dct_8x8_stage_2_0_t428 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t442;
    FSM_dct_8x8_stage_2_0_t444 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_2_0_t445 = FSM_dct_8x8_stage_2_0_t444[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t446 = FSM_dct_8x8_stage_2_0_t445 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_2_0_t447 = FSM_dct_8x8_stage_2_0_t446[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t448 = FSM_dct_8x8_stage_2_0_t447[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t449 = FSM_dct_8x8_stage_2_0_t443;
    FSM_dct_8x8_stage_2_0_t449[FSM_dct_8x8_stage_2_0_t448 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t434 - FSM_dct_8x8_stage_2_0_t440;
    FSM_dct_8x8_stage_2_0_t450 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_2_0_t451 = FSM_dct_8x8_stage_2_0_t450[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t452 = FSM_dct_8x8_stage_2_0_t451 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_2_0_t453 = FSM_dct_8x8_stage_2_0_t452[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t454 = FSM_dct_8x8_stage_2_0_t453[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t455 = FSM_dct_8x8_stage_2_0_t449;
    FSM_dct_8x8_stage_2_0_t455[FSM_dct_8x8_stage_2_0_t454 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t414 - FSM_dct_8x8_stage_2_0_t420;
    FSM_dct_8x8_stage_2_0_t456 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_2_0_t457 = FSM_dct_8x8_stage_2_0_t456[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t458 = FSM_dct_8x8_stage_2_0_t457 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_2_0_t459 = FSM_dct_8x8_stage_2_0_t458[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t460 = FSM_dct_8x8_stage_2_0_t459[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t461 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_2_0_t462 = FSM_dct_8x8_stage_2_0_t461[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t463 = FSM_dct_8x8_stage_2_0_t462 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_2_0_t464 = FSM_dct_8x8_stage_2_0_t463[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t465 = FSM_dct_8x8_stage_2_0_t464[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t466 = i_data_in[FSM_dct_8x8_stage_2_0_t465 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t467 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_2_0_t468 = FSM_dct_8x8_stage_2_0_t467[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t469 = FSM_dct_8x8_stage_2_0_t468 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_2_0_t470 = FSM_dct_8x8_stage_2_0_t469[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t471 = FSM_dct_8x8_stage_2_0_t470[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t472 = i_data_in[FSM_dct_8x8_stage_2_0_t471 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t473 = FSM_dct_8x8_stage_2_0_t466 + FSM_dct_8x8_stage_2_0_t472;
    FSM_dct_8x8_stage_2_0_t474 = FSM_dct_8x8_stage_2_0_t473[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t475 = FSM_dct_8x8_stage_2_0_t455;
    FSM_dct_8x8_stage_2_0_t475[FSM_dct_8x8_stage_2_0_t460 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t474;
    FSM_dct_8x8_stage_2_0_t476 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_2_0_t477 = FSM_dct_8x8_stage_2_0_t476[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t478 = FSM_dct_8x8_stage_2_0_t477 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_2_0_t479 = FSM_dct_8x8_stage_2_0_t478[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t480 = FSM_dct_8x8_stage_2_0_t479[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t481 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_2_0_t482 = FSM_dct_8x8_stage_2_0_t481[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t483 = FSM_dct_8x8_stage_2_0_t482 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_2_0_t484 = FSM_dct_8x8_stage_2_0_t483[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t485 = FSM_dct_8x8_stage_2_0_t484[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t486 = i_data_in[FSM_dct_8x8_stage_2_0_t485 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t487 = FSM_dct_8x8_stage_2_0_t472 + FSM_dct_8x8_stage_2_0_t486;
    FSM_dct_8x8_stage_2_0_t488 = FSM_dct_8x8_stage_2_0_t487[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t489 = FSM_dct_8x8_stage_2_0_t475;
    FSM_dct_8x8_stage_2_0_t489[FSM_dct_8x8_stage_2_0_t480 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t488;
    FSM_dct_8x8_stage_2_0_t490 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_2_0_t491 = FSM_dct_8x8_stage_2_0_t490[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t492 = FSM_dct_8x8_stage_2_0_t491 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_2_0_t493 = FSM_dct_8x8_stage_2_0_t492[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t494 = FSM_dct_8x8_stage_2_0_t493[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t495 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_2_0_t496 = FSM_dct_8x8_stage_2_0_t495[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t497 = FSM_dct_8x8_stage_2_0_t496 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_2_0_t498 = FSM_dct_8x8_stage_2_0_t497[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t499 = FSM_dct_8x8_stage_2_0_t498[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t500 = i_data_in[FSM_dct_8x8_stage_2_0_t499 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t501 = FSM_dct_8x8_stage_2_0_t486 + FSM_dct_8x8_stage_2_0_t500;
    FSM_dct_8x8_stage_2_0_t502 = FSM_dct_8x8_stage_2_0_t501[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t503 = FSM_dct_8x8_stage_2_0_t489;
    FSM_dct_8x8_stage_2_0_t503[FSM_dct_8x8_stage_2_0_t494 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t502;
    FSM_dct_8x8_stage_2_0_t504 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_2_0_t505 = FSM_dct_8x8_stage_2_0_t504[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t506 = FSM_dct_8x8_stage_2_0_t505 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_2_0_t507 = FSM_dct_8x8_stage_2_0_t506[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t508 = FSM_dct_8x8_stage_2_0_t507[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t509 = FSM_dct_8x8_stage_2_0_t503;
    FSM_dct_8x8_stage_2_0_t509[FSM_dct_8x8_stage_2_0_t508 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t500;
    FSM_dct_8x8_stage_2_0_t510 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_2_0_t511 = FSM_dct_8x8_stage_2_0_t510[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t512 = FSM_dct_8x8_stage_2_0_t511[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t513 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_2_0_t514 = FSM_dct_8x8_stage_2_0_t513[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t515 = FSM_dct_8x8_stage_2_0_t514[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t516 = i_data_in[FSM_dct_8x8_stage_2_0_t515 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t517 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_2_0_t518 = FSM_dct_8x8_stage_2_0_t517[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t519 = FSM_dct_8x8_stage_2_0_t518 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_2_0_t520 = FSM_dct_8x8_stage_2_0_t519[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t521 = FSM_dct_8x8_stage_2_0_t520[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t522 = i_data_in[FSM_dct_8x8_stage_2_0_t521 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t523 = FSM_dct_8x8_stage_2_0_t516 + FSM_dct_8x8_stage_2_0_t522;
    FSM_dct_8x8_stage_2_0_t524 = FSM_dct_8x8_stage_2_0_t523[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t525 = FSM_dct_8x8_stage_2_0_t509;
    FSM_dct_8x8_stage_2_0_t525[FSM_dct_8x8_stage_2_0_t512 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t524;
    FSM_dct_8x8_stage_2_0_t526 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_2_0_t527 = FSM_dct_8x8_stage_2_0_t526[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t528 = FSM_dct_8x8_stage_2_0_t527 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_2_0_t529 = FSM_dct_8x8_stage_2_0_t528[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t530 = FSM_dct_8x8_stage_2_0_t529[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t531 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_2_0_t532 = FSM_dct_8x8_stage_2_0_t531[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t533 = FSM_dct_8x8_stage_2_0_t532 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_2_0_t534 = FSM_dct_8x8_stage_2_0_t533[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t535 = FSM_dct_8x8_stage_2_0_t534[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t536 = i_data_in[FSM_dct_8x8_stage_2_0_t535 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t537 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_2_0_t538 = FSM_dct_8x8_stage_2_0_t537[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t539 = FSM_dct_8x8_stage_2_0_t538 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_2_0_t540 = FSM_dct_8x8_stage_2_0_t539[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t541 = FSM_dct_8x8_stage_2_0_t540[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t542 = i_data_in[FSM_dct_8x8_stage_2_0_t541 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t543 = FSM_dct_8x8_stage_2_0_t536 + FSM_dct_8x8_stage_2_0_t542;
    FSM_dct_8x8_stage_2_0_t544 = FSM_dct_8x8_stage_2_0_t543[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t545 = FSM_dct_8x8_stage_2_0_t525;
    FSM_dct_8x8_stage_2_0_t545[FSM_dct_8x8_stage_2_0_t530 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t544;
    FSM_dct_8x8_stage_2_0_t546 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_2_0_t547 = FSM_dct_8x8_stage_2_0_t546[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t548 = FSM_dct_8x8_stage_2_0_t547 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_2_0_t549 = FSM_dct_8x8_stage_2_0_t548[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t550 = FSM_dct_8x8_stage_2_0_t549[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t551 = FSM_dct_8x8_stage_2_0_t545;
    FSM_dct_8x8_stage_2_0_t551[FSM_dct_8x8_stage_2_0_t550 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t536 - FSM_dct_8x8_stage_2_0_t542;
    FSM_dct_8x8_stage_2_0_t552 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_2_0_t553 = FSM_dct_8x8_stage_2_0_t552[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t554 = FSM_dct_8x8_stage_2_0_t553 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_2_0_t555 = FSM_dct_8x8_stage_2_0_t554[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t556 = FSM_dct_8x8_stage_2_0_t555[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t557 = FSM_dct_8x8_stage_2_0_t551;
    FSM_dct_8x8_stage_2_0_t557[FSM_dct_8x8_stage_2_0_t556 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t516 - FSM_dct_8x8_stage_2_0_t522;
    FSM_dct_8x8_stage_2_0_t558 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_2_0_t559 = FSM_dct_8x8_stage_2_0_t558[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t560 = FSM_dct_8x8_stage_2_0_t559 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_2_0_t561 = FSM_dct_8x8_stage_2_0_t560[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t562 = FSM_dct_8x8_stage_2_0_t561[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t563 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_2_0_t564 = FSM_dct_8x8_stage_2_0_t563[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t565 = FSM_dct_8x8_stage_2_0_t564 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_2_0_t566 = FSM_dct_8x8_stage_2_0_t565[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t567 = FSM_dct_8x8_stage_2_0_t566[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t568 = i_data_in[FSM_dct_8x8_stage_2_0_t567 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t569 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_2_0_t570 = FSM_dct_8x8_stage_2_0_t569[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t571 = FSM_dct_8x8_stage_2_0_t570 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_2_0_t572 = FSM_dct_8x8_stage_2_0_t571[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t573 = FSM_dct_8x8_stage_2_0_t572[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t574 = i_data_in[FSM_dct_8x8_stage_2_0_t573 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t575 = FSM_dct_8x8_stage_2_0_t568 + FSM_dct_8x8_stage_2_0_t574;
    FSM_dct_8x8_stage_2_0_t576 = FSM_dct_8x8_stage_2_0_t575[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t577 = FSM_dct_8x8_stage_2_0_t557;
    FSM_dct_8x8_stage_2_0_t577[FSM_dct_8x8_stage_2_0_t562 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t576;
    FSM_dct_8x8_stage_2_0_t578 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_2_0_t579 = FSM_dct_8x8_stage_2_0_t578[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t580 = FSM_dct_8x8_stage_2_0_t579 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_2_0_t581 = FSM_dct_8x8_stage_2_0_t580[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t582 = FSM_dct_8x8_stage_2_0_t581[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t583 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_2_0_t584 = FSM_dct_8x8_stage_2_0_t583[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t585 = FSM_dct_8x8_stage_2_0_t584 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_2_0_t586 = FSM_dct_8x8_stage_2_0_t585[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t587 = FSM_dct_8x8_stage_2_0_t586[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t588 = i_data_in[FSM_dct_8x8_stage_2_0_t587 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t589 = FSM_dct_8x8_stage_2_0_t574 + FSM_dct_8x8_stage_2_0_t588;
    FSM_dct_8x8_stage_2_0_t590 = FSM_dct_8x8_stage_2_0_t589[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t591 = FSM_dct_8x8_stage_2_0_t577;
    FSM_dct_8x8_stage_2_0_t591[FSM_dct_8x8_stage_2_0_t582 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t590;
    FSM_dct_8x8_stage_2_0_t592 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_2_0_t593 = FSM_dct_8x8_stage_2_0_t592[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t594 = FSM_dct_8x8_stage_2_0_t593 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_2_0_t595 = FSM_dct_8x8_stage_2_0_t594[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t596 = FSM_dct_8x8_stage_2_0_t595[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t597 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_2_0_t598 = FSM_dct_8x8_stage_2_0_t597[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t599 = FSM_dct_8x8_stage_2_0_t598 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_2_0_t600 = FSM_dct_8x8_stage_2_0_t599[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t601 = FSM_dct_8x8_stage_2_0_t600[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t602 = i_data_in[FSM_dct_8x8_stage_2_0_t601 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t603 = FSM_dct_8x8_stage_2_0_t588 + FSM_dct_8x8_stage_2_0_t602;
    FSM_dct_8x8_stage_2_0_t604 = FSM_dct_8x8_stage_2_0_t603[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t605 = FSM_dct_8x8_stage_2_0_t591;
    FSM_dct_8x8_stage_2_0_t605[FSM_dct_8x8_stage_2_0_t596 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t604;
    FSM_dct_8x8_stage_2_0_t606 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_2_0_t607 = FSM_dct_8x8_stage_2_0_t606[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t608 = FSM_dct_8x8_stage_2_0_t607 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_2_0_t609 = FSM_dct_8x8_stage_2_0_t608[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t610 = FSM_dct_8x8_stage_2_0_t609[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t611 = FSM_dct_8x8_stage_2_0_t605;
    FSM_dct_8x8_stage_2_0_t611[FSM_dct_8x8_stage_2_0_t610 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t602;
    FSM_dct_8x8_stage_2_0_t612 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_2_0_t613 = FSM_dct_8x8_stage_2_0_t612[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t614 = FSM_dct_8x8_stage_2_0_t613[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t615 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_2_0_t616 = FSM_dct_8x8_stage_2_0_t615[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t617 = FSM_dct_8x8_stage_2_0_t616[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t618 = i_data_in[FSM_dct_8x8_stage_2_0_t617 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t619 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_2_0_t620 = FSM_dct_8x8_stage_2_0_t619[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t621 = FSM_dct_8x8_stage_2_0_t620 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_2_0_t622 = FSM_dct_8x8_stage_2_0_t621[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t623 = FSM_dct_8x8_stage_2_0_t622[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t624 = i_data_in[FSM_dct_8x8_stage_2_0_t623 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t625 = FSM_dct_8x8_stage_2_0_t618 + FSM_dct_8x8_stage_2_0_t624;
    FSM_dct_8x8_stage_2_0_t626 = FSM_dct_8x8_stage_2_0_t625[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t627 = FSM_dct_8x8_stage_2_0_t611;
    FSM_dct_8x8_stage_2_0_t627[FSM_dct_8x8_stage_2_0_t614 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t626;
    FSM_dct_8x8_stage_2_0_t628 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_2_0_t629 = FSM_dct_8x8_stage_2_0_t628[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t630 = FSM_dct_8x8_stage_2_0_t629 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_2_0_t631 = FSM_dct_8x8_stage_2_0_t630[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t632 = FSM_dct_8x8_stage_2_0_t631[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t633 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_2_0_t634 = FSM_dct_8x8_stage_2_0_t633[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t635 = FSM_dct_8x8_stage_2_0_t634 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_2_0_t636 = FSM_dct_8x8_stage_2_0_t635[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t637 = FSM_dct_8x8_stage_2_0_t636[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t638 = i_data_in[FSM_dct_8x8_stage_2_0_t637 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t639 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_2_0_t640 = FSM_dct_8x8_stage_2_0_t639[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t641 = FSM_dct_8x8_stage_2_0_t640 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_2_0_t642 = FSM_dct_8x8_stage_2_0_t641[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t643 = FSM_dct_8x8_stage_2_0_t642[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t644 = i_data_in[FSM_dct_8x8_stage_2_0_t643 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t645 = FSM_dct_8x8_stage_2_0_t638 + FSM_dct_8x8_stage_2_0_t644;
    FSM_dct_8x8_stage_2_0_t646 = FSM_dct_8x8_stage_2_0_t645[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t647 = FSM_dct_8x8_stage_2_0_t627;
    FSM_dct_8x8_stage_2_0_t647[FSM_dct_8x8_stage_2_0_t632 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t646;
    FSM_dct_8x8_stage_2_0_t648 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_2_0_t649 = FSM_dct_8x8_stage_2_0_t648[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t650 = FSM_dct_8x8_stage_2_0_t649 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_2_0_t651 = FSM_dct_8x8_stage_2_0_t650[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t652 = FSM_dct_8x8_stage_2_0_t651[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t653 = FSM_dct_8x8_stage_2_0_t647;
    FSM_dct_8x8_stage_2_0_t653[FSM_dct_8x8_stage_2_0_t652 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t638 - FSM_dct_8x8_stage_2_0_t644;
    FSM_dct_8x8_stage_2_0_t654 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_2_0_t655 = FSM_dct_8x8_stage_2_0_t654[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t656 = FSM_dct_8x8_stage_2_0_t655 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_2_0_t657 = FSM_dct_8x8_stage_2_0_t656[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t658 = FSM_dct_8x8_stage_2_0_t657[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t659 = FSM_dct_8x8_stage_2_0_t653;
    FSM_dct_8x8_stage_2_0_t659[FSM_dct_8x8_stage_2_0_t658 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t618 - FSM_dct_8x8_stage_2_0_t624;
    FSM_dct_8x8_stage_2_0_t660 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_2_0_t661 = FSM_dct_8x8_stage_2_0_t660[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t662 = FSM_dct_8x8_stage_2_0_t661 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_2_0_t663 = FSM_dct_8x8_stage_2_0_t662[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t664 = FSM_dct_8x8_stage_2_0_t663[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t665 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_2_0_t666 = FSM_dct_8x8_stage_2_0_t665[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t667 = FSM_dct_8x8_stage_2_0_t666 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_2_0_t668 = FSM_dct_8x8_stage_2_0_t667[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t669 = FSM_dct_8x8_stage_2_0_t668[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t670 = i_data_in[FSM_dct_8x8_stage_2_0_t669 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t671 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_2_0_t672 = FSM_dct_8x8_stage_2_0_t671[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t673 = FSM_dct_8x8_stage_2_0_t672 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_2_0_t674 = FSM_dct_8x8_stage_2_0_t673[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t675 = FSM_dct_8x8_stage_2_0_t674[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t676 = i_data_in[FSM_dct_8x8_stage_2_0_t675 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t677 = FSM_dct_8x8_stage_2_0_t670 + FSM_dct_8x8_stage_2_0_t676;
    FSM_dct_8x8_stage_2_0_t678 = FSM_dct_8x8_stage_2_0_t677[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t679 = FSM_dct_8x8_stage_2_0_t659;
    FSM_dct_8x8_stage_2_0_t679[FSM_dct_8x8_stage_2_0_t664 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t678;
    FSM_dct_8x8_stage_2_0_t680 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_2_0_t681 = FSM_dct_8x8_stage_2_0_t680[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t682 = FSM_dct_8x8_stage_2_0_t681 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_2_0_t683 = FSM_dct_8x8_stage_2_0_t682[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t684 = FSM_dct_8x8_stage_2_0_t683[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t685 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_2_0_t686 = FSM_dct_8x8_stage_2_0_t685[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t687 = FSM_dct_8x8_stage_2_0_t686 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_2_0_t688 = FSM_dct_8x8_stage_2_0_t687[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t689 = FSM_dct_8x8_stage_2_0_t688[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t690 = i_data_in[FSM_dct_8x8_stage_2_0_t689 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t691 = FSM_dct_8x8_stage_2_0_t676 + FSM_dct_8x8_stage_2_0_t690;
    FSM_dct_8x8_stage_2_0_t692 = FSM_dct_8x8_stage_2_0_t691[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t693 = FSM_dct_8x8_stage_2_0_t679;
    FSM_dct_8x8_stage_2_0_t693[FSM_dct_8x8_stage_2_0_t684 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t692;
    FSM_dct_8x8_stage_2_0_t694 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_2_0_t695 = FSM_dct_8x8_stage_2_0_t694[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t696 = FSM_dct_8x8_stage_2_0_t695 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_2_0_t697 = FSM_dct_8x8_stage_2_0_t696[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t698 = FSM_dct_8x8_stage_2_0_t697[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t699 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_2_0_t700 = FSM_dct_8x8_stage_2_0_t699[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t701 = FSM_dct_8x8_stage_2_0_t700 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_2_0_t702 = FSM_dct_8x8_stage_2_0_t701[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t703 = FSM_dct_8x8_stage_2_0_t702[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t704 = i_data_in[FSM_dct_8x8_stage_2_0_t703 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t705 = FSM_dct_8x8_stage_2_0_t690 + FSM_dct_8x8_stage_2_0_t704;
    FSM_dct_8x8_stage_2_0_t706 = FSM_dct_8x8_stage_2_0_t705[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t707 = FSM_dct_8x8_stage_2_0_t693;
    FSM_dct_8x8_stage_2_0_t707[FSM_dct_8x8_stage_2_0_t698 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t706;
    FSM_dct_8x8_stage_2_0_t708 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_2_0_t709 = FSM_dct_8x8_stage_2_0_t708[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t710 = FSM_dct_8x8_stage_2_0_t709 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_2_0_t711 = FSM_dct_8x8_stage_2_0_t710[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t712 = FSM_dct_8x8_stage_2_0_t711[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t713 = FSM_dct_8x8_stage_2_0_t707;
    FSM_dct_8x8_stage_2_0_t713[FSM_dct_8x8_stage_2_0_t712 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t704;
    FSM_dct_8x8_stage_2_0_t714 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_2_0_t715 = FSM_dct_8x8_stage_2_0_t714[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t716 = FSM_dct_8x8_stage_2_0_t715[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t717 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_2_0_t718 = FSM_dct_8x8_stage_2_0_t717[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t719 = FSM_dct_8x8_stage_2_0_t718[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t720 = i_data_in[FSM_dct_8x8_stage_2_0_t719 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t721 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_2_0_t722 = FSM_dct_8x8_stage_2_0_t721[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t723 = FSM_dct_8x8_stage_2_0_t722 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_2_0_t724 = FSM_dct_8x8_stage_2_0_t723[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t725 = FSM_dct_8x8_stage_2_0_t724[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t726 = i_data_in[FSM_dct_8x8_stage_2_0_t725 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t727 = FSM_dct_8x8_stage_2_0_t720 + FSM_dct_8x8_stage_2_0_t726;
    FSM_dct_8x8_stage_2_0_t728 = FSM_dct_8x8_stage_2_0_t727[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t729 = FSM_dct_8x8_stage_2_0_t713;
    FSM_dct_8x8_stage_2_0_t729[FSM_dct_8x8_stage_2_0_t716 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t728;
    FSM_dct_8x8_stage_2_0_t730 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_2_0_t731 = FSM_dct_8x8_stage_2_0_t730[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t732 = FSM_dct_8x8_stage_2_0_t731 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_2_0_t733 = FSM_dct_8x8_stage_2_0_t732[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t734 = FSM_dct_8x8_stage_2_0_t733[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t735 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_2_0_t736 = FSM_dct_8x8_stage_2_0_t735[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t737 = FSM_dct_8x8_stage_2_0_t736 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_2_0_t738 = FSM_dct_8x8_stage_2_0_t737[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t739 = FSM_dct_8x8_stage_2_0_t738[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t740 = i_data_in[FSM_dct_8x8_stage_2_0_t739 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t741 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_2_0_t742 = FSM_dct_8x8_stage_2_0_t741[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t743 = FSM_dct_8x8_stage_2_0_t742 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_2_0_t744 = FSM_dct_8x8_stage_2_0_t743[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t745 = FSM_dct_8x8_stage_2_0_t744[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t746 = i_data_in[FSM_dct_8x8_stage_2_0_t745 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t747 = FSM_dct_8x8_stage_2_0_t740 + FSM_dct_8x8_stage_2_0_t746;
    FSM_dct_8x8_stage_2_0_t748 = FSM_dct_8x8_stage_2_0_t747[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t749 = FSM_dct_8x8_stage_2_0_t729;
    FSM_dct_8x8_stage_2_0_t749[FSM_dct_8x8_stage_2_0_t734 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t748;
    FSM_dct_8x8_stage_2_0_t750 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_2_0_t751 = FSM_dct_8x8_stage_2_0_t750[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t752 = FSM_dct_8x8_stage_2_0_t751 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_2_0_t753 = FSM_dct_8x8_stage_2_0_t752[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t754 = FSM_dct_8x8_stage_2_0_t753[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t755 = FSM_dct_8x8_stage_2_0_t749;
    FSM_dct_8x8_stage_2_0_t755[FSM_dct_8x8_stage_2_0_t754 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t740 - FSM_dct_8x8_stage_2_0_t746;
    FSM_dct_8x8_stage_2_0_t756 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_2_0_t757 = FSM_dct_8x8_stage_2_0_t756[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t758 = FSM_dct_8x8_stage_2_0_t757 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_2_0_t759 = FSM_dct_8x8_stage_2_0_t758[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t760 = FSM_dct_8x8_stage_2_0_t759[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t761 = FSM_dct_8x8_stage_2_0_t755;
    FSM_dct_8x8_stage_2_0_t761[FSM_dct_8x8_stage_2_0_t760 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t720 - FSM_dct_8x8_stage_2_0_t726;
    FSM_dct_8x8_stage_2_0_t762 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_2_0_t763 = FSM_dct_8x8_stage_2_0_t762[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t764 = FSM_dct_8x8_stage_2_0_t763 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_2_0_t765 = FSM_dct_8x8_stage_2_0_t764[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t766 = FSM_dct_8x8_stage_2_0_t765[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t767 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_2_0_t768 = FSM_dct_8x8_stage_2_0_t767[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t769 = FSM_dct_8x8_stage_2_0_t768 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_2_0_t770 = FSM_dct_8x8_stage_2_0_t769[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t771 = FSM_dct_8x8_stage_2_0_t770[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t772 = i_data_in[FSM_dct_8x8_stage_2_0_t771 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t773 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_2_0_t774 = FSM_dct_8x8_stage_2_0_t773[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t775 = FSM_dct_8x8_stage_2_0_t774 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_2_0_t776 = FSM_dct_8x8_stage_2_0_t775[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t777 = FSM_dct_8x8_stage_2_0_t776[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t778 = i_data_in[FSM_dct_8x8_stage_2_0_t777 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t779 = FSM_dct_8x8_stage_2_0_t772 + FSM_dct_8x8_stage_2_0_t778;
    FSM_dct_8x8_stage_2_0_t780 = FSM_dct_8x8_stage_2_0_t779[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t781 = FSM_dct_8x8_stage_2_0_t761;
    FSM_dct_8x8_stage_2_0_t781[FSM_dct_8x8_stage_2_0_t766 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t780;
    FSM_dct_8x8_stage_2_0_t782 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_2_0_t783 = FSM_dct_8x8_stage_2_0_t782[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t784 = FSM_dct_8x8_stage_2_0_t783 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_2_0_t785 = FSM_dct_8x8_stage_2_0_t784[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t786 = FSM_dct_8x8_stage_2_0_t785[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t787 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_2_0_t788 = FSM_dct_8x8_stage_2_0_t787[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t789 = FSM_dct_8x8_stage_2_0_t788 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_2_0_t790 = FSM_dct_8x8_stage_2_0_t789[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t791 = FSM_dct_8x8_stage_2_0_t790[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t792 = i_data_in[FSM_dct_8x8_stage_2_0_t791 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t793 = FSM_dct_8x8_stage_2_0_t778 + FSM_dct_8x8_stage_2_0_t792;
    FSM_dct_8x8_stage_2_0_t794 = FSM_dct_8x8_stage_2_0_t793[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t795 = FSM_dct_8x8_stage_2_0_t781;
    FSM_dct_8x8_stage_2_0_t795[FSM_dct_8x8_stage_2_0_t786 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t794;
    FSM_dct_8x8_stage_2_0_t796 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_2_0_t797 = FSM_dct_8x8_stage_2_0_t796[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t798 = FSM_dct_8x8_stage_2_0_t797 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_2_0_t799 = FSM_dct_8x8_stage_2_0_t798[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t800 = FSM_dct_8x8_stage_2_0_t799[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t801 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_2_0_t802 = FSM_dct_8x8_stage_2_0_t801[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t803 = FSM_dct_8x8_stage_2_0_t802 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_2_0_t804 = FSM_dct_8x8_stage_2_0_t803[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t805 = FSM_dct_8x8_stage_2_0_t804[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t806 = i_data_in[FSM_dct_8x8_stage_2_0_t805 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t807 = FSM_dct_8x8_stage_2_0_t792 + FSM_dct_8x8_stage_2_0_t806;
    FSM_dct_8x8_stage_2_0_t808 = FSM_dct_8x8_stage_2_0_t807[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t809 = FSM_dct_8x8_stage_2_0_t795;
    FSM_dct_8x8_stage_2_0_t809[FSM_dct_8x8_stage_2_0_t800 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t808;
    FSM_dct_8x8_stage_2_0_t810 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_2_0_t811 = FSM_dct_8x8_stage_2_0_t810[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t812 = FSM_dct_8x8_stage_2_0_t811 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_2_0_t813 = FSM_dct_8x8_stage_2_0_t812[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t814 = FSM_dct_8x8_stage_2_0_t813[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t815 = FSM_dct_8x8_stage_2_0_t809;
    FSM_dct_8x8_stage_2_0_t815[FSM_dct_8x8_stage_2_0_t814 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t806;
end

always @* begin
    FSM_dct_8x8_stage_2_0_t0 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_2_0_t1 = FSM_dct_8x8_stage_2_0_t0[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t2 = FSM_dct_8x8_stage_2_0_t1[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t3 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_2_0_t4 = FSM_dct_8x8_stage_2_0_t3[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t5 = FSM_dct_8x8_stage_2_0_t4[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t6 = i_data_in[FSM_dct_8x8_stage_2_0_t5 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t7 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_2_0_t8 = FSM_dct_8x8_stage_2_0_t7[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t9 = FSM_dct_8x8_stage_2_0_t8 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_2_0_t10 = FSM_dct_8x8_stage_2_0_t9[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t11 = FSM_dct_8x8_stage_2_0_t10[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t12 = i_data_in[FSM_dct_8x8_stage_2_0_t11 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t13 = FSM_dct_8x8_stage_2_0_t6 + FSM_dct_8x8_stage_2_0_t12;
    FSM_dct_8x8_stage_2_0_t14 = FSM_dct_8x8_stage_2_0_t13[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t15 = 2048'b0;
    FSM_dct_8x8_stage_2_0_t15[FSM_dct_8x8_stage_2_0_t2 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t14;
    FSM_dct_8x8_stage_2_0_t16 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_2_0_t17 = FSM_dct_8x8_stage_2_0_t16[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t18 = FSM_dct_8x8_stage_2_0_t17 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_2_0_t19 = FSM_dct_8x8_stage_2_0_t18[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t20 = FSM_dct_8x8_stage_2_0_t19[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t21 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_2_0_t22 = FSM_dct_8x8_stage_2_0_t21[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t23 = FSM_dct_8x8_stage_2_0_t22 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_2_0_t24 = FSM_dct_8x8_stage_2_0_t23[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t25 = FSM_dct_8x8_stage_2_0_t24[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t26 = i_data_in[FSM_dct_8x8_stage_2_0_t25 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t27 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_2_0_t28 = FSM_dct_8x8_stage_2_0_t27[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t29 = FSM_dct_8x8_stage_2_0_t28 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_2_0_t30 = FSM_dct_8x8_stage_2_0_t29[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t31 = FSM_dct_8x8_stage_2_0_t30[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t32 = i_data_in[FSM_dct_8x8_stage_2_0_t31 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t33 = FSM_dct_8x8_stage_2_0_t26 + FSM_dct_8x8_stage_2_0_t32;
    FSM_dct_8x8_stage_2_0_t34 = FSM_dct_8x8_stage_2_0_t33[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t35 = FSM_dct_8x8_stage_2_0_t15;
    FSM_dct_8x8_stage_2_0_t35[FSM_dct_8x8_stage_2_0_t20 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t34;
    FSM_dct_8x8_stage_2_0_t36 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_2_0_t37 = FSM_dct_8x8_stage_2_0_t36[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t38 = FSM_dct_8x8_stage_2_0_t37 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_2_0_t39 = FSM_dct_8x8_stage_2_0_t38[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t40 = FSM_dct_8x8_stage_2_0_t39[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t41 = FSM_dct_8x8_stage_2_0_t35;
    FSM_dct_8x8_stage_2_0_t41[FSM_dct_8x8_stage_2_0_t40 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t26 - FSM_dct_8x8_stage_2_0_t32;
    FSM_dct_8x8_stage_2_0_t42 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_2_0_t43 = FSM_dct_8x8_stage_2_0_t42[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t44 = FSM_dct_8x8_stage_2_0_t43 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_2_0_t45 = FSM_dct_8x8_stage_2_0_t44[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t46 = FSM_dct_8x8_stage_2_0_t45[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t47 = FSM_dct_8x8_stage_2_0_t41;
    FSM_dct_8x8_stage_2_0_t47[FSM_dct_8x8_stage_2_0_t46 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t6 - FSM_dct_8x8_stage_2_0_t12;
    FSM_dct_8x8_stage_2_0_t48 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_2_0_t49 = FSM_dct_8x8_stage_2_0_t48[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t50 = FSM_dct_8x8_stage_2_0_t49 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_2_0_t51 = FSM_dct_8x8_stage_2_0_t50[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t52 = FSM_dct_8x8_stage_2_0_t51[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t53 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_2_0_t54 = FSM_dct_8x8_stage_2_0_t53[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t55 = FSM_dct_8x8_stage_2_0_t54 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_2_0_t56 = FSM_dct_8x8_stage_2_0_t55[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t57 = FSM_dct_8x8_stage_2_0_t56[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t58 = i_data_in[FSM_dct_8x8_stage_2_0_t57 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t59 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_2_0_t60 = FSM_dct_8x8_stage_2_0_t59[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t61 = FSM_dct_8x8_stage_2_0_t60 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_2_0_t62 = FSM_dct_8x8_stage_2_0_t61[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t63 = FSM_dct_8x8_stage_2_0_t62[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t64 = i_data_in[FSM_dct_8x8_stage_2_0_t63 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t65 = FSM_dct_8x8_stage_2_0_t58 + FSM_dct_8x8_stage_2_0_t64;
    FSM_dct_8x8_stage_2_0_t66 = FSM_dct_8x8_stage_2_0_t65[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t67 = FSM_dct_8x8_stage_2_0_t47;
    FSM_dct_8x8_stage_2_0_t67[FSM_dct_8x8_stage_2_0_t52 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t66;
    FSM_dct_8x8_stage_2_0_t68 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_2_0_t69 = FSM_dct_8x8_stage_2_0_t68[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t70 = FSM_dct_8x8_stage_2_0_t69 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_2_0_t71 = FSM_dct_8x8_stage_2_0_t70[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t72 = FSM_dct_8x8_stage_2_0_t71[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t73 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_2_0_t74 = FSM_dct_8x8_stage_2_0_t73[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t75 = FSM_dct_8x8_stage_2_0_t74 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_2_0_t76 = FSM_dct_8x8_stage_2_0_t75[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t77 = FSM_dct_8x8_stage_2_0_t76[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t78 = i_data_in[FSM_dct_8x8_stage_2_0_t77 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t79 = FSM_dct_8x8_stage_2_0_t64 + FSM_dct_8x8_stage_2_0_t78;
    FSM_dct_8x8_stage_2_0_t80 = FSM_dct_8x8_stage_2_0_t79[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t81 = FSM_dct_8x8_stage_2_0_t67;
    FSM_dct_8x8_stage_2_0_t81[FSM_dct_8x8_stage_2_0_t72 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t80;
    FSM_dct_8x8_stage_2_0_t82 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_2_0_t83 = FSM_dct_8x8_stage_2_0_t82[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t84 = FSM_dct_8x8_stage_2_0_t83 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_2_0_t85 = FSM_dct_8x8_stage_2_0_t84[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t86 = FSM_dct_8x8_stage_2_0_t85[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t87 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_2_0_t88 = FSM_dct_8x8_stage_2_0_t87[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t89 = FSM_dct_8x8_stage_2_0_t88 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_2_0_t90 = FSM_dct_8x8_stage_2_0_t89[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t91 = FSM_dct_8x8_stage_2_0_t90[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t92 = i_data_in[FSM_dct_8x8_stage_2_0_t91 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t93 = FSM_dct_8x8_stage_2_0_t78 + FSM_dct_8x8_stage_2_0_t92;
    FSM_dct_8x8_stage_2_0_t94 = FSM_dct_8x8_stage_2_0_t93[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t95 = FSM_dct_8x8_stage_2_0_t81;
    FSM_dct_8x8_stage_2_0_t95[FSM_dct_8x8_stage_2_0_t86 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t94;
    FSM_dct_8x8_stage_2_0_t96 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_2_0_t97 = FSM_dct_8x8_stage_2_0_t96[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t98 = FSM_dct_8x8_stage_2_0_t97 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_2_0_t99 = FSM_dct_8x8_stage_2_0_t98[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t100 = FSM_dct_8x8_stage_2_0_t99[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t101 = FSM_dct_8x8_stage_2_0_t95;
    FSM_dct_8x8_stage_2_0_t101[FSM_dct_8x8_stage_2_0_t100 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t92;
    FSM_dct_8x8_stage_2_0_t102 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_2_0_t103 = FSM_dct_8x8_stage_2_0_t102[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t104 = FSM_dct_8x8_stage_2_0_t103[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t105 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_2_0_t106 = FSM_dct_8x8_stage_2_0_t105[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t107 = FSM_dct_8x8_stage_2_0_t106[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t108 = i_data_in[FSM_dct_8x8_stage_2_0_t107 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t109 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_2_0_t110 = FSM_dct_8x8_stage_2_0_t109[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t111 = FSM_dct_8x8_stage_2_0_t110 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_2_0_t112 = FSM_dct_8x8_stage_2_0_t111[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t113 = FSM_dct_8x8_stage_2_0_t112[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t114 = i_data_in[FSM_dct_8x8_stage_2_0_t113 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t115 = FSM_dct_8x8_stage_2_0_t108 + FSM_dct_8x8_stage_2_0_t114;
    FSM_dct_8x8_stage_2_0_t116 = FSM_dct_8x8_stage_2_0_t115[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t117 = FSM_dct_8x8_stage_2_0_t101;
    FSM_dct_8x8_stage_2_0_t117[FSM_dct_8x8_stage_2_0_t104 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t116;
    FSM_dct_8x8_stage_2_0_t118 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_2_0_t119 = FSM_dct_8x8_stage_2_0_t118[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t120 = FSM_dct_8x8_stage_2_0_t119 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_2_0_t121 = FSM_dct_8x8_stage_2_0_t120[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t122 = FSM_dct_8x8_stage_2_0_t121[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t123 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_2_0_t124 = FSM_dct_8x8_stage_2_0_t123[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t125 = FSM_dct_8x8_stage_2_0_t124 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_2_0_t126 = FSM_dct_8x8_stage_2_0_t125[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t127 = FSM_dct_8x8_stage_2_0_t126[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t128 = i_data_in[FSM_dct_8x8_stage_2_0_t127 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t129 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_2_0_t130 = FSM_dct_8x8_stage_2_0_t129[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t131 = FSM_dct_8x8_stage_2_0_t130 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_2_0_t132 = FSM_dct_8x8_stage_2_0_t131[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t133 = FSM_dct_8x8_stage_2_0_t132[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t134 = i_data_in[FSM_dct_8x8_stage_2_0_t133 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t135 = FSM_dct_8x8_stage_2_0_t128 + FSM_dct_8x8_stage_2_0_t134;
    FSM_dct_8x8_stage_2_0_t136 = FSM_dct_8x8_stage_2_0_t135[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t137 = FSM_dct_8x8_stage_2_0_t117;
    FSM_dct_8x8_stage_2_0_t137[FSM_dct_8x8_stage_2_0_t122 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t136;
    FSM_dct_8x8_stage_2_0_t138 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_2_0_t139 = FSM_dct_8x8_stage_2_0_t138[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t140 = FSM_dct_8x8_stage_2_0_t139 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_2_0_t141 = FSM_dct_8x8_stage_2_0_t140[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t142 = FSM_dct_8x8_stage_2_0_t141[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t143 = FSM_dct_8x8_stage_2_0_t137;
    FSM_dct_8x8_stage_2_0_t143[FSM_dct_8x8_stage_2_0_t142 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t128 - FSM_dct_8x8_stage_2_0_t134;
    FSM_dct_8x8_stage_2_0_t144 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_2_0_t145 = FSM_dct_8x8_stage_2_0_t144[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t146 = FSM_dct_8x8_stage_2_0_t145 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_2_0_t147 = FSM_dct_8x8_stage_2_0_t146[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t148 = FSM_dct_8x8_stage_2_0_t147[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t149 = FSM_dct_8x8_stage_2_0_t143;
    FSM_dct_8x8_stage_2_0_t149[FSM_dct_8x8_stage_2_0_t148 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t108 - FSM_dct_8x8_stage_2_0_t114;
    FSM_dct_8x8_stage_2_0_t150 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_2_0_t151 = FSM_dct_8x8_stage_2_0_t150[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t152 = FSM_dct_8x8_stage_2_0_t151 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_2_0_t153 = FSM_dct_8x8_stage_2_0_t152[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t154 = FSM_dct_8x8_stage_2_0_t153[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t155 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_2_0_t156 = FSM_dct_8x8_stage_2_0_t155[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t157 = FSM_dct_8x8_stage_2_0_t156 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_2_0_t158 = FSM_dct_8x8_stage_2_0_t157[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t159 = FSM_dct_8x8_stage_2_0_t158[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t160 = i_data_in[FSM_dct_8x8_stage_2_0_t159 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t161 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_2_0_t162 = FSM_dct_8x8_stage_2_0_t161[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t163 = FSM_dct_8x8_stage_2_0_t162 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_2_0_t164 = FSM_dct_8x8_stage_2_0_t163[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t165 = FSM_dct_8x8_stage_2_0_t164[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t166 = i_data_in[FSM_dct_8x8_stage_2_0_t165 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t167 = FSM_dct_8x8_stage_2_0_t160 + FSM_dct_8x8_stage_2_0_t166;
    FSM_dct_8x8_stage_2_0_t168 = FSM_dct_8x8_stage_2_0_t167[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t169 = FSM_dct_8x8_stage_2_0_t149;
    FSM_dct_8x8_stage_2_0_t169[FSM_dct_8x8_stage_2_0_t154 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t168;
    FSM_dct_8x8_stage_2_0_t170 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_2_0_t171 = FSM_dct_8x8_stage_2_0_t170[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t172 = FSM_dct_8x8_stage_2_0_t171 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_2_0_t173 = FSM_dct_8x8_stage_2_0_t172[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t174 = FSM_dct_8x8_stage_2_0_t173[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t175 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_2_0_t176 = FSM_dct_8x8_stage_2_0_t175[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t177 = FSM_dct_8x8_stage_2_0_t176 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_2_0_t178 = FSM_dct_8x8_stage_2_0_t177[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t179 = FSM_dct_8x8_stage_2_0_t178[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t180 = i_data_in[FSM_dct_8x8_stage_2_0_t179 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t181 = FSM_dct_8x8_stage_2_0_t166 + FSM_dct_8x8_stage_2_0_t180;
    FSM_dct_8x8_stage_2_0_t182 = FSM_dct_8x8_stage_2_0_t181[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t183 = FSM_dct_8x8_stage_2_0_t169;
    FSM_dct_8x8_stage_2_0_t183[FSM_dct_8x8_stage_2_0_t174 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t182;
    FSM_dct_8x8_stage_2_0_t184 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_2_0_t185 = FSM_dct_8x8_stage_2_0_t184[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t186 = FSM_dct_8x8_stage_2_0_t185 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_2_0_t187 = FSM_dct_8x8_stage_2_0_t186[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t188 = FSM_dct_8x8_stage_2_0_t187[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t189 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_2_0_t190 = FSM_dct_8x8_stage_2_0_t189[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t191 = FSM_dct_8x8_stage_2_0_t190 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_2_0_t192 = FSM_dct_8x8_stage_2_0_t191[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t193 = FSM_dct_8x8_stage_2_0_t192[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t194 = i_data_in[FSM_dct_8x8_stage_2_0_t193 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t195 = FSM_dct_8x8_stage_2_0_t180 + FSM_dct_8x8_stage_2_0_t194;
    FSM_dct_8x8_stage_2_0_t196 = FSM_dct_8x8_stage_2_0_t195[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t197 = FSM_dct_8x8_stage_2_0_t183;
    FSM_dct_8x8_stage_2_0_t197[FSM_dct_8x8_stage_2_0_t188 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t196;
    FSM_dct_8x8_stage_2_0_t198 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_2_0_t199 = FSM_dct_8x8_stage_2_0_t198[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t200 = FSM_dct_8x8_stage_2_0_t199 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_2_0_t201 = FSM_dct_8x8_stage_2_0_t200[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t202 = FSM_dct_8x8_stage_2_0_t201[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t203 = FSM_dct_8x8_stage_2_0_t197;
    FSM_dct_8x8_stage_2_0_t203[FSM_dct_8x8_stage_2_0_t202 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t194;
    FSM_dct_8x8_stage_2_0_t204 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_2_0_t205 = FSM_dct_8x8_stage_2_0_t204[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t206 = FSM_dct_8x8_stage_2_0_t205[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t207 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_2_0_t208 = FSM_dct_8x8_stage_2_0_t207[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t209 = FSM_dct_8x8_stage_2_0_t208[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t210 = i_data_in[FSM_dct_8x8_stage_2_0_t209 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t211 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_2_0_t212 = FSM_dct_8x8_stage_2_0_t211[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t213 = FSM_dct_8x8_stage_2_0_t212 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_2_0_t214 = FSM_dct_8x8_stage_2_0_t213[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t215 = FSM_dct_8x8_stage_2_0_t214[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t216 = i_data_in[FSM_dct_8x8_stage_2_0_t215 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t217 = FSM_dct_8x8_stage_2_0_t210 + FSM_dct_8x8_stage_2_0_t216;
    FSM_dct_8x8_stage_2_0_t218 = FSM_dct_8x8_stage_2_0_t217[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t219 = FSM_dct_8x8_stage_2_0_t203;
    FSM_dct_8x8_stage_2_0_t219[FSM_dct_8x8_stage_2_0_t206 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t218;
    FSM_dct_8x8_stage_2_0_t220 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_2_0_t221 = FSM_dct_8x8_stage_2_0_t220[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t222 = FSM_dct_8x8_stage_2_0_t221 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_2_0_t223 = FSM_dct_8x8_stage_2_0_t222[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t224 = FSM_dct_8x8_stage_2_0_t223[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t225 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_2_0_t226 = FSM_dct_8x8_stage_2_0_t225[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t227 = FSM_dct_8x8_stage_2_0_t226 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_2_0_t228 = FSM_dct_8x8_stage_2_0_t227[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t229 = FSM_dct_8x8_stage_2_0_t228[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t230 = i_data_in[FSM_dct_8x8_stage_2_0_t229 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t231 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_2_0_t232 = FSM_dct_8x8_stage_2_0_t231[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t233 = FSM_dct_8x8_stage_2_0_t232 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_2_0_t234 = FSM_dct_8x8_stage_2_0_t233[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t235 = FSM_dct_8x8_stage_2_0_t234[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t236 = i_data_in[FSM_dct_8x8_stage_2_0_t235 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t237 = FSM_dct_8x8_stage_2_0_t230 + FSM_dct_8x8_stage_2_0_t236;
    FSM_dct_8x8_stage_2_0_t238 = FSM_dct_8x8_stage_2_0_t237[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t239 = FSM_dct_8x8_stage_2_0_t219;
    FSM_dct_8x8_stage_2_0_t239[FSM_dct_8x8_stage_2_0_t224 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t238;
    FSM_dct_8x8_stage_2_0_t240 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_2_0_t241 = FSM_dct_8x8_stage_2_0_t240[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t242 = FSM_dct_8x8_stage_2_0_t241 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_2_0_t243 = FSM_dct_8x8_stage_2_0_t242[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t244 = FSM_dct_8x8_stage_2_0_t243[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t245 = FSM_dct_8x8_stage_2_0_t239;
    FSM_dct_8x8_stage_2_0_t245[FSM_dct_8x8_stage_2_0_t244 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t230 - FSM_dct_8x8_stage_2_0_t236;
    FSM_dct_8x8_stage_2_0_t246 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_2_0_t247 = FSM_dct_8x8_stage_2_0_t246[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t248 = FSM_dct_8x8_stage_2_0_t247 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_2_0_t249 = FSM_dct_8x8_stage_2_0_t248[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t250 = FSM_dct_8x8_stage_2_0_t249[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t251 = FSM_dct_8x8_stage_2_0_t245;
    FSM_dct_8x8_stage_2_0_t251[FSM_dct_8x8_stage_2_0_t250 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t210 - FSM_dct_8x8_stage_2_0_t216;
    FSM_dct_8x8_stage_2_0_t252 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_2_0_t253 = FSM_dct_8x8_stage_2_0_t252[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t254 = FSM_dct_8x8_stage_2_0_t253 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_2_0_t255 = FSM_dct_8x8_stage_2_0_t254[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t256 = FSM_dct_8x8_stage_2_0_t255[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t257 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_2_0_t258 = FSM_dct_8x8_stage_2_0_t257[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t259 = FSM_dct_8x8_stage_2_0_t258 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_2_0_t260 = FSM_dct_8x8_stage_2_0_t259[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t261 = FSM_dct_8x8_stage_2_0_t260[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t262 = i_data_in[FSM_dct_8x8_stage_2_0_t261 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t263 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_2_0_t264 = FSM_dct_8x8_stage_2_0_t263[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t265 = FSM_dct_8x8_stage_2_0_t264 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_2_0_t266 = FSM_dct_8x8_stage_2_0_t265[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t267 = FSM_dct_8x8_stage_2_0_t266[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t268 = i_data_in[FSM_dct_8x8_stage_2_0_t267 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t269 = FSM_dct_8x8_stage_2_0_t262 + FSM_dct_8x8_stage_2_0_t268;
    FSM_dct_8x8_stage_2_0_t270 = FSM_dct_8x8_stage_2_0_t269[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t271 = FSM_dct_8x8_stage_2_0_t251;
    FSM_dct_8x8_stage_2_0_t271[FSM_dct_8x8_stage_2_0_t256 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t270;
    FSM_dct_8x8_stage_2_0_t272 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_2_0_t273 = FSM_dct_8x8_stage_2_0_t272[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t274 = FSM_dct_8x8_stage_2_0_t273 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_2_0_t275 = FSM_dct_8x8_stage_2_0_t274[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t276 = FSM_dct_8x8_stage_2_0_t275[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t277 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_2_0_t278 = FSM_dct_8x8_stage_2_0_t277[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t279 = FSM_dct_8x8_stage_2_0_t278 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_2_0_t280 = FSM_dct_8x8_stage_2_0_t279[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t281 = FSM_dct_8x8_stage_2_0_t280[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t282 = i_data_in[FSM_dct_8x8_stage_2_0_t281 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t283 = FSM_dct_8x8_stage_2_0_t268 + FSM_dct_8x8_stage_2_0_t282;
    FSM_dct_8x8_stage_2_0_t284 = FSM_dct_8x8_stage_2_0_t283[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t285 = FSM_dct_8x8_stage_2_0_t271;
    FSM_dct_8x8_stage_2_0_t285[FSM_dct_8x8_stage_2_0_t276 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t284;
    FSM_dct_8x8_stage_2_0_t286 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_2_0_t287 = FSM_dct_8x8_stage_2_0_t286[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t288 = FSM_dct_8x8_stage_2_0_t287 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_2_0_t289 = FSM_dct_8x8_stage_2_0_t288[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t290 = FSM_dct_8x8_stage_2_0_t289[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t291 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_2_0_t292 = FSM_dct_8x8_stage_2_0_t291[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t293 = FSM_dct_8x8_stage_2_0_t292 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_2_0_t294 = FSM_dct_8x8_stage_2_0_t293[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t295 = FSM_dct_8x8_stage_2_0_t294[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t296 = i_data_in[FSM_dct_8x8_stage_2_0_t295 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t297 = FSM_dct_8x8_stage_2_0_t282 + FSM_dct_8x8_stage_2_0_t296;
    FSM_dct_8x8_stage_2_0_t298 = FSM_dct_8x8_stage_2_0_t297[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t299 = FSM_dct_8x8_stage_2_0_t285;
    FSM_dct_8x8_stage_2_0_t299[FSM_dct_8x8_stage_2_0_t290 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t298;
    FSM_dct_8x8_stage_2_0_t300 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_2_0_t301 = FSM_dct_8x8_stage_2_0_t300[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t302 = FSM_dct_8x8_stage_2_0_t301 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_2_0_t303 = FSM_dct_8x8_stage_2_0_t302[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t304 = FSM_dct_8x8_stage_2_0_t303[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t305 = FSM_dct_8x8_stage_2_0_t299;
    FSM_dct_8x8_stage_2_0_t305[FSM_dct_8x8_stage_2_0_t304 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t296;
    FSM_dct_8x8_stage_2_0_t306 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_2_0_t307 = FSM_dct_8x8_stage_2_0_t306[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t308 = FSM_dct_8x8_stage_2_0_t307[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t309 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_2_0_t310 = FSM_dct_8x8_stage_2_0_t309[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t311 = FSM_dct_8x8_stage_2_0_t310[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t312 = i_data_in[FSM_dct_8x8_stage_2_0_t311 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t313 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_2_0_t314 = FSM_dct_8x8_stage_2_0_t313[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t315 = FSM_dct_8x8_stage_2_0_t314 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_2_0_t316 = FSM_dct_8x8_stage_2_0_t315[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t317 = FSM_dct_8x8_stage_2_0_t316[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t318 = i_data_in[FSM_dct_8x8_stage_2_0_t317 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t319 = FSM_dct_8x8_stage_2_0_t312 + FSM_dct_8x8_stage_2_0_t318;
    FSM_dct_8x8_stage_2_0_t320 = FSM_dct_8x8_stage_2_0_t319[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t321 = FSM_dct_8x8_stage_2_0_t305;
    FSM_dct_8x8_stage_2_0_t321[FSM_dct_8x8_stage_2_0_t308 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t320;
    FSM_dct_8x8_stage_2_0_t322 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_2_0_t323 = FSM_dct_8x8_stage_2_0_t322[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t324 = FSM_dct_8x8_stage_2_0_t323 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_2_0_t325 = FSM_dct_8x8_stage_2_0_t324[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t326 = FSM_dct_8x8_stage_2_0_t325[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t327 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_2_0_t328 = FSM_dct_8x8_stage_2_0_t327[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t329 = FSM_dct_8x8_stage_2_0_t328 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_2_0_t330 = FSM_dct_8x8_stage_2_0_t329[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t331 = FSM_dct_8x8_stage_2_0_t330[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t332 = i_data_in[FSM_dct_8x8_stage_2_0_t331 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t333 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_2_0_t334 = FSM_dct_8x8_stage_2_0_t333[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t335 = FSM_dct_8x8_stage_2_0_t334 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_2_0_t336 = FSM_dct_8x8_stage_2_0_t335[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t337 = FSM_dct_8x8_stage_2_0_t336[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t338 = i_data_in[FSM_dct_8x8_stage_2_0_t337 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t339 = FSM_dct_8x8_stage_2_0_t332 + FSM_dct_8x8_stage_2_0_t338;
    FSM_dct_8x8_stage_2_0_t340 = FSM_dct_8x8_stage_2_0_t339[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t341 = FSM_dct_8x8_stage_2_0_t321;
    FSM_dct_8x8_stage_2_0_t341[FSM_dct_8x8_stage_2_0_t326 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t340;
    FSM_dct_8x8_stage_2_0_t342 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_2_0_t343 = FSM_dct_8x8_stage_2_0_t342[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t344 = FSM_dct_8x8_stage_2_0_t343 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_2_0_t345 = FSM_dct_8x8_stage_2_0_t344[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t346 = FSM_dct_8x8_stage_2_0_t345[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t347 = FSM_dct_8x8_stage_2_0_t341;
    FSM_dct_8x8_stage_2_0_t347[FSM_dct_8x8_stage_2_0_t346 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t332 - FSM_dct_8x8_stage_2_0_t338;
    FSM_dct_8x8_stage_2_0_t348 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_2_0_t349 = FSM_dct_8x8_stage_2_0_t348[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t350 = FSM_dct_8x8_stage_2_0_t349 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_2_0_t351 = FSM_dct_8x8_stage_2_0_t350[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t352 = FSM_dct_8x8_stage_2_0_t351[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t353 = FSM_dct_8x8_stage_2_0_t347;
    FSM_dct_8x8_stage_2_0_t353[FSM_dct_8x8_stage_2_0_t352 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t312 - FSM_dct_8x8_stage_2_0_t318;
    FSM_dct_8x8_stage_2_0_t354 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_2_0_t355 = FSM_dct_8x8_stage_2_0_t354[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t356 = FSM_dct_8x8_stage_2_0_t355 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_2_0_t357 = FSM_dct_8x8_stage_2_0_t356[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t358 = FSM_dct_8x8_stage_2_0_t357[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t359 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_2_0_t360 = FSM_dct_8x8_stage_2_0_t359[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t361 = FSM_dct_8x8_stage_2_0_t360 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_2_0_t362 = FSM_dct_8x8_stage_2_0_t361[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t363 = FSM_dct_8x8_stage_2_0_t362[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t364 = i_data_in[FSM_dct_8x8_stage_2_0_t363 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t365 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_2_0_t366 = FSM_dct_8x8_stage_2_0_t365[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t367 = FSM_dct_8x8_stage_2_0_t366 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_2_0_t368 = FSM_dct_8x8_stage_2_0_t367[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t369 = FSM_dct_8x8_stage_2_0_t368[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t370 = i_data_in[FSM_dct_8x8_stage_2_0_t369 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t371 = FSM_dct_8x8_stage_2_0_t364 + FSM_dct_8x8_stage_2_0_t370;
    FSM_dct_8x8_stage_2_0_t372 = FSM_dct_8x8_stage_2_0_t371[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t373 = FSM_dct_8x8_stage_2_0_t353;
    FSM_dct_8x8_stage_2_0_t373[FSM_dct_8x8_stage_2_0_t358 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t372;
    FSM_dct_8x8_stage_2_0_t374 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_2_0_t375 = FSM_dct_8x8_stage_2_0_t374[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t376 = FSM_dct_8x8_stage_2_0_t375 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_2_0_t377 = FSM_dct_8x8_stage_2_0_t376[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t378 = FSM_dct_8x8_stage_2_0_t377[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t379 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_2_0_t380 = FSM_dct_8x8_stage_2_0_t379[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t381 = FSM_dct_8x8_stage_2_0_t380 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_2_0_t382 = FSM_dct_8x8_stage_2_0_t381[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t383 = FSM_dct_8x8_stage_2_0_t382[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t384 = i_data_in[FSM_dct_8x8_stage_2_0_t383 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t385 = FSM_dct_8x8_stage_2_0_t370 + FSM_dct_8x8_stage_2_0_t384;
    FSM_dct_8x8_stage_2_0_t386 = FSM_dct_8x8_stage_2_0_t385[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t387 = FSM_dct_8x8_stage_2_0_t373;
    FSM_dct_8x8_stage_2_0_t387[FSM_dct_8x8_stage_2_0_t378 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t386;
    FSM_dct_8x8_stage_2_0_t388 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_2_0_t389 = FSM_dct_8x8_stage_2_0_t388[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t390 = FSM_dct_8x8_stage_2_0_t389 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_2_0_t391 = FSM_dct_8x8_stage_2_0_t390[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t392 = FSM_dct_8x8_stage_2_0_t391[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t393 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_2_0_t394 = FSM_dct_8x8_stage_2_0_t393[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t395 = FSM_dct_8x8_stage_2_0_t394 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_2_0_t396 = FSM_dct_8x8_stage_2_0_t395[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t397 = FSM_dct_8x8_stage_2_0_t396[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t398 = i_data_in[FSM_dct_8x8_stage_2_0_t397 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t399 = FSM_dct_8x8_stage_2_0_t384 + FSM_dct_8x8_stage_2_0_t398;
    FSM_dct_8x8_stage_2_0_t400 = FSM_dct_8x8_stage_2_0_t399[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t401 = FSM_dct_8x8_stage_2_0_t387;
    FSM_dct_8x8_stage_2_0_t401[FSM_dct_8x8_stage_2_0_t392 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t400;
    FSM_dct_8x8_stage_2_0_t402 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_2_0_t403 = FSM_dct_8x8_stage_2_0_t402[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t404 = FSM_dct_8x8_stage_2_0_t403 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_2_0_t405 = FSM_dct_8x8_stage_2_0_t404[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t406 = FSM_dct_8x8_stage_2_0_t405[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t407 = FSM_dct_8x8_stage_2_0_t401;
    FSM_dct_8x8_stage_2_0_t407[FSM_dct_8x8_stage_2_0_t406 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t398;
    FSM_dct_8x8_stage_2_0_t408 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_2_0_t409 = FSM_dct_8x8_stage_2_0_t408[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t410 = FSM_dct_8x8_stage_2_0_t409[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t411 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_2_0_t412 = FSM_dct_8x8_stage_2_0_t411[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t413 = FSM_dct_8x8_stage_2_0_t412[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t414 = i_data_in[FSM_dct_8x8_stage_2_0_t413 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t415 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_2_0_t416 = FSM_dct_8x8_stage_2_0_t415[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t417 = FSM_dct_8x8_stage_2_0_t416 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_2_0_t418 = FSM_dct_8x8_stage_2_0_t417[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t419 = FSM_dct_8x8_stage_2_0_t418[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t420 = i_data_in[FSM_dct_8x8_stage_2_0_t419 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t421 = FSM_dct_8x8_stage_2_0_t414 + FSM_dct_8x8_stage_2_0_t420;
    FSM_dct_8x8_stage_2_0_t422 = FSM_dct_8x8_stage_2_0_t421[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t423 = FSM_dct_8x8_stage_2_0_t407;
    FSM_dct_8x8_stage_2_0_t423[FSM_dct_8x8_stage_2_0_t410 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t422;
    FSM_dct_8x8_stage_2_0_t424 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_2_0_t425 = FSM_dct_8x8_stage_2_0_t424[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t426 = FSM_dct_8x8_stage_2_0_t425 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_2_0_t427 = FSM_dct_8x8_stage_2_0_t426[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t428 = FSM_dct_8x8_stage_2_0_t427[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t429 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_2_0_t430 = FSM_dct_8x8_stage_2_0_t429[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t431 = FSM_dct_8x8_stage_2_0_t430 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_2_0_t432 = FSM_dct_8x8_stage_2_0_t431[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t433 = FSM_dct_8x8_stage_2_0_t432[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t434 = i_data_in[FSM_dct_8x8_stage_2_0_t433 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t435 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_2_0_t436 = FSM_dct_8x8_stage_2_0_t435[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t437 = FSM_dct_8x8_stage_2_0_t436 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_2_0_t438 = FSM_dct_8x8_stage_2_0_t437[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t439 = FSM_dct_8x8_stage_2_0_t438[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t440 = i_data_in[FSM_dct_8x8_stage_2_0_t439 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t441 = FSM_dct_8x8_stage_2_0_t434 + FSM_dct_8x8_stage_2_0_t440;
    FSM_dct_8x8_stage_2_0_t442 = FSM_dct_8x8_stage_2_0_t441[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t443 = FSM_dct_8x8_stage_2_0_t423;
    FSM_dct_8x8_stage_2_0_t443[FSM_dct_8x8_stage_2_0_t428 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t442;
    FSM_dct_8x8_stage_2_0_t444 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_2_0_t445 = FSM_dct_8x8_stage_2_0_t444[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t446 = FSM_dct_8x8_stage_2_0_t445 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_2_0_t447 = FSM_dct_8x8_stage_2_0_t446[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t448 = FSM_dct_8x8_stage_2_0_t447[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t449 = FSM_dct_8x8_stage_2_0_t443;
    FSM_dct_8x8_stage_2_0_t449[FSM_dct_8x8_stage_2_0_t448 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t434 - FSM_dct_8x8_stage_2_0_t440;
    FSM_dct_8x8_stage_2_0_t450 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_2_0_t451 = FSM_dct_8x8_stage_2_0_t450[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t452 = FSM_dct_8x8_stage_2_0_t451 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_2_0_t453 = FSM_dct_8x8_stage_2_0_t452[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t454 = FSM_dct_8x8_stage_2_0_t453[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t455 = FSM_dct_8x8_stage_2_0_t449;
    FSM_dct_8x8_stage_2_0_t455[FSM_dct_8x8_stage_2_0_t454 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t414 - FSM_dct_8x8_stage_2_0_t420;
    FSM_dct_8x8_stage_2_0_t456 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_2_0_t457 = FSM_dct_8x8_stage_2_0_t456[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t458 = FSM_dct_8x8_stage_2_0_t457 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_2_0_t459 = FSM_dct_8x8_stage_2_0_t458[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t460 = FSM_dct_8x8_stage_2_0_t459[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t461 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_2_0_t462 = FSM_dct_8x8_stage_2_0_t461[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t463 = FSM_dct_8x8_stage_2_0_t462 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_2_0_t464 = FSM_dct_8x8_stage_2_0_t463[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t465 = FSM_dct_8x8_stage_2_0_t464[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t466 = i_data_in[FSM_dct_8x8_stage_2_0_t465 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t467 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_2_0_t468 = FSM_dct_8x8_stage_2_0_t467[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t469 = FSM_dct_8x8_stage_2_0_t468 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_2_0_t470 = FSM_dct_8x8_stage_2_0_t469[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t471 = FSM_dct_8x8_stage_2_0_t470[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t472 = i_data_in[FSM_dct_8x8_stage_2_0_t471 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t473 = FSM_dct_8x8_stage_2_0_t466 + FSM_dct_8x8_stage_2_0_t472;
    FSM_dct_8x8_stage_2_0_t474 = FSM_dct_8x8_stage_2_0_t473[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t475 = FSM_dct_8x8_stage_2_0_t455;
    FSM_dct_8x8_stage_2_0_t475[FSM_dct_8x8_stage_2_0_t460 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t474;
    FSM_dct_8x8_stage_2_0_t476 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_2_0_t477 = FSM_dct_8x8_stage_2_0_t476[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t478 = FSM_dct_8x8_stage_2_0_t477 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_2_0_t479 = FSM_dct_8x8_stage_2_0_t478[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t480 = FSM_dct_8x8_stage_2_0_t479[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t481 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_2_0_t482 = FSM_dct_8x8_stage_2_0_t481[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t483 = FSM_dct_8x8_stage_2_0_t482 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_2_0_t484 = FSM_dct_8x8_stage_2_0_t483[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t485 = FSM_dct_8x8_stage_2_0_t484[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t486 = i_data_in[FSM_dct_8x8_stage_2_0_t485 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t487 = FSM_dct_8x8_stage_2_0_t472 + FSM_dct_8x8_stage_2_0_t486;
    FSM_dct_8x8_stage_2_0_t488 = FSM_dct_8x8_stage_2_0_t487[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t489 = FSM_dct_8x8_stage_2_0_t475;
    FSM_dct_8x8_stage_2_0_t489[FSM_dct_8x8_stage_2_0_t480 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t488;
    FSM_dct_8x8_stage_2_0_t490 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_2_0_t491 = FSM_dct_8x8_stage_2_0_t490[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t492 = FSM_dct_8x8_stage_2_0_t491 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_2_0_t493 = FSM_dct_8x8_stage_2_0_t492[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t494 = FSM_dct_8x8_stage_2_0_t493[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t495 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_2_0_t496 = FSM_dct_8x8_stage_2_0_t495[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t497 = FSM_dct_8x8_stage_2_0_t496 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_2_0_t498 = FSM_dct_8x8_stage_2_0_t497[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t499 = FSM_dct_8x8_stage_2_0_t498[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t500 = i_data_in[FSM_dct_8x8_stage_2_0_t499 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t501 = FSM_dct_8x8_stage_2_0_t486 + FSM_dct_8x8_stage_2_0_t500;
    FSM_dct_8x8_stage_2_0_t502 = FSM_dct_8x8_stage_2_0_t501[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t503 = FSM_dct_8x8_stage_2_0_t489;
    FSM_dct_8x8_stage_2_0_t503[FSM_dct_8x8_stage_2_0_t494 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t502;
    FSM_dct_8x8_stage_2_0_t504 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_2_0_t505 = FSM_dct_8x8_stage_2_0_t504[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t506 = FSM_dct_8x8_stage_2_0_t505 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_2_0_t507 = FSM_dct_8x8_stage_2_0_t506[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t508 = FSM_dct_8x8_stage_2_0_t507[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t509 = FSM_dct_8x8_stage_2_0_t503;
    FSM_dct_8x8_stage_2_0_t509[FSM_dct_8x8_stage_2_0_t508 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t500;
    FSM_dct_8x8_stage_2_0_t510 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_2_0_t511 = FSM_dct_8x8_stage_2_0_t510[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t512 = FSM_dct_8x8_stage_2_0_t511[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t513 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_2_0_t514 = FSM_dct_8x8_stage_2_0_t513[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t515 = FSM_dct_8x8_stage_2_0_t514[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t516 = i_data_in[FSM_dct_8x8_stage_2_0_t515 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t517 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_2_0_t518 = FSM_dct_8x8_stage_2_0_t517[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t519 = FSM_dct_8x8_stage_2_0_t518 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_2_0_t520 = FSM_dct_8x8_stage_2_0_t519[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t521 = FSM_dct_8x8_stage_2_0_t520[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t522 = i_data_in[FSM_dct_8x8_stage_2_0_t521 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t523 = FSM_dct_8x8_stage_2_0_t516 + FSM_dct_8x8_stage_2_0_t522;
    FSM_dct_8x8_stage_2_0_t524 = FSM_dct_8x8_stage_2_0_t523[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t525 = FSM_dct_8x8_stage_2_0_t509;
    FSM_dct_8x8_stage_2_0_t525[FSM_dct_8x8_stage_2_0_t512 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t524;
    FSM_dct_8x8_stage_2_0_t526 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_2_0_t527 = FSM_dct_8x8_stage_2_0_t526[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t528 = FSM_dct_8x8_stage_2_0_t527 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_2_0_t529 = FSM_dct_8x8_stage_2_0_t528[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t530 = FSM_dct_8x8_stage_2_0_t529[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t531 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_2_0_t532 = FSM_dct_8x8_stage_2_0_t531[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t533 = FSM_dct_8x8_stage_2_0_t532 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_2_0_t534 = FSM_dct_8x8_stage_2_0_t533[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t535 = FSM_dct_8x8_stage_2_0_t534[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t536 = i_data_in[FSM_dct_8x8_stage_2_0_t535 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t537 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_2_0_t538 = FSM_dct_8x8_stage_2_0_t537[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t539 = FSM_dct_8x8_stage_2_0_t538 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_2_0_t540 = FSM_dct_8x8_stage_2_0_t539[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t541 = FSM_dct_8x8_stage_2_0_t540[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t542 = i_data_in[FSM_dct_8x8_stage_2_0_t541 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t543 = FSM_dct_8x8_stage_2_0_t536 + FSM_dct_8x8_stage_2_0_t542;
    FSM_dct_8x8_stage_2_0_t544 = FSM_dct_8x8_stage_2_0_t543[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t545 = FSM_dct_8x8_stage_2_0_t525;
    FSM_dct_8x8_stage_2_0_t545[FSM_dct_8x8_stage_2_0_t530 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t544;
    FSM_dct_8x8_stage_2_0_t546 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_2_0_t547 = FSM_dct_8x8_stage_2_0_t546[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t548 = FSM_dct_8x8_stage_2_0_t547 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_2_0_t549 = FSM_dct_8x8_stage_2_0_t548[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t550 = FSM_dct_8x8_stage_2_0_t549[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t551 = FSM_dct_8x8_stage_2_0_t545;
    FSM_dct_8x8_stage_2_0_t551[FSM_dct_8x8_stage_2_0_t550 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t536 - FSM_dct_8x8_stage_2_0_t542;
    FSM_dct_8x8_stage_2_0_t552 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_2_0_t553 = FSM_dct_8x8_stage_2_0_t552[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t554 = FSM_dct_8x8_stage_2_0_t553 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_2_0_t555 = FSM_dct_8x8_stage_2_0_t554[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t556 = FSM_dct_8x8_stage_2_0_t555[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t557 = FSM_dct_8x8_stage_2_0_t551;
    FSM_dct_8x8_stage_2_0_t557[FSM_dct_8x8_stage_2_0_t556 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t516 - FSM_dct_8x8_stage_2_0_t522;
    FSM_dct_8x8_stage_2_0_t558 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_2_0_t559 = FSM_dct_8x8_stage_2_0_t558[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t560 = FSM_dct_8x8_stage_2_0_t559 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_2_0_t561 = FSM_dct_8x8_stage_2_0_t560[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t562 = FSM_dct_8x8_stage_2_0_t561[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t563 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_2_0_t564 = FSM_dct_8x8_stage_2_0_t563[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t565 = FSM_dct_8x8_stage_2_0_t564 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_2_0_t566 = FSM_dct_8x8_stage_2_0_t565[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t567 = FSM_dct_8x8_stage_2_0_t566[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t568 = i_data_in[FSM_dct_8x8_stage_2_0_t567 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t569 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_2_0_t570 = FSM_dct_8x8_stage_2_0_t569[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t571 = FSM_dct_8x8_stage_2_0_t570 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_2_0_t572 = FSM_dct_8x8_stage_2_0_t571[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t573 = FSM_dct_8x8_stage_2_0_t572[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t574 = i_data_in[FSM_dct_8x8_stage_2_0_t573 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t575 = FSM_dct_8x8_stage_2_0_t568 + FSM_dct_8x8_stage_2_0_t574;
    FSM_dct_8x8_stage_2_0_t576 = FSM_dct_8x8_stage_2_0_t575[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t577 = FSM_dct_8x8_stage_2_0_t557;
    FSM_dct_8x8_stage_2_0_t577[FSM_dct_8x8_stage_2_0_t562 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t576;
    FSM_dct_8x8_stage_2_0_t578 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_2_0_t579 = FSM_dct_8x8_stage_2_0_t578[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t580 = FSM_dct_8x8_stage_2_0_t579 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_2_0_t581 = FSM_dct_8x8_stage_2_0_t580[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t582 = FSM_dct_8x8_stage_2_0_t581[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t583 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_2_0_t584 = FSM_dct_8x8_stage_2_0_t583[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t585 = FSM_dct_8x8_stage_2_0_t584 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_2_0_t586 = FSM_dct_8x8_stage_2_0_t585[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t587 = FSM_dct_8x8_stage_2_0_t586[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t588 = i_data_in[FSM_dct_8x8_stage_2_0_t587 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t589 = FSM_dct_8x8_stage_2_0_t574 + FSM_dct_8x8_stage_2_0_t588;
    FSM_dct_8x8_stage_2_0_t590 = FSM_dct_8x8_stage_2_0_t589[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t591 = FSM_dct_8x8_stage_2_0_t577;
    FSM_dct_8x8_stage_2_0_t591[FSM_dct_8x8_stage_2_0_t582 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t590;
    FSM_dct_8x8_stage_2_0_t592 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_2_0_t593 = FSM_dct_8x8_stage_2_0_t592[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t594 = FSM_dct_8x8_stage_2_0_t593 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_2_0_t595 = FSM_dct_8x8_stage_2_0_t594[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t596 = FSM_dct_8x8_stage_2_0_t595[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t597 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_2_0_t598 = FSM_dct_8x8_stage_2_0_t597[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t599 = FSM_dct_8x8_stage_2_0_t598 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_2_0_t600 = FSM_dct_8x8_stage_2_0_t599[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t601 = FSM_dct_8x8_stage_2_0_t600[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t602 = i_data_in[FSM_dct_8x8_stage_2_0_t601 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t603 = FSM_dct_8x8_stage_2_0_t588 + FSM_dct_8x8_stage_2_0_t602;
    FSM_dct_8x8_stage_2_0_t604 = FSM_dct_8x8_stage_2_0_t603[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t605 = FSM_dct_8x8_stage_2_0_t591;
    FSM_dct_8x8_stage_2_0_t605[FSM_dct_8x8_stage_2_0_t596 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t604;
    FSM_dct_8x8_stage_2_0_t606 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_2_0_t607 = FSM_dct_8x8_stage_2_0_t606[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t608 = FSM_dct_8x8_stage_2_0_t607 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_2_0_t609 = FSM_dct_8x8_stage_2_0_t608[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t610 = FSM_dct_8x8_stage_2_0_t609[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t611 = FSM_dct_8x8_stage_2_0_t605;
    FSM_dct_8x8_stage_2_0_t611[FSM_dct_8x8_stage_2_0_t610 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t602;
    FSM_dct_8x8_stage_2_0_t612 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_2_0_t613 = FSM_dct_8x8_stage_2_0_t612[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t614 = FSM_dct_8x8_stage_2_0_t613[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t615 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_2_0_t616 = FSM_dct_8x8_stage_2_0_t615[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t617 = FSM_dct_8x8_stage_2_0_t616[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t618 = i_data_in[FSM_dct_8x8_stage_2_0_t617 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t619 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_2_0_t620 = FSM_dct_8x8_stage_2_0_t619[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t621 = FSM_dct_8x8_stage_2_0_t620 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_2_0_t622 = FSM_dct_8x8_stage_2_0_t621[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t623 = FSM_dct_8x8_stage_2_0_t622[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t624 = i_data_in[FSM_dct_8x8_stage_2_0_t623 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t625 = FSM_dct_8x8_stage_2_0_t618 + FSM_dct_8x8_stage_2_0_t624;
    FSM_dct_8x8_stage_2_0_t626 = FSM_dct_8x8_stage_2_0_t625[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t627 = FSM_dct_8x8_stage_2_0_t611;
    FSM_dct_8x8_stage_2_0_t627[FSM_dct_8x8_stage_2_0_t614 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t626;
    FSM_dct_8x8_stage_2_0_t628 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_2_0_t629 = FSM_dct_8x8_stage_2_0_t628[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t630 = FSM_dct_8x8_stage_2_0_t629 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_2_0_t631 = FSM_dct_8x8_stage_2_0_t630[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t632 = FSM_dct_8x8_stage_2_0_t631[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t633 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_2_0_t634 = FSM_dct_8x8_stage_2_0_t633[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t635 = FSM_dct_8x8_stage_2_0_t634 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_2_0_t636 = FSM_dct_8x8_stage_2_0_t635[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t637 = FSM_dct_8x8_stage_2_0_t636[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t638 = i_data_in[FSM_dct_8x8_stage_2_0_t637 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t639 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_2_0_t640 = FSM_dct_8x8_stage_2_0_t639[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t641 = FSM_dct_8x8_stage_2_0_t640 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_2_0_t642 = FSM_dct_8x8_stage_2_0_t641[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t643 = FSM_dct_8x8_stage_2_0_t642[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t644 = i_data_in[FSM_dct_8x8_stage_2_0_t643 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t645 = FSM_dct_8x8_stage_2_0_t638 + FSM_dct_8x8_stage_2_0_t644;
    FSM_dct_8x8_stage_2_0_t646 = FSM_dct_8x8_stage_2_0_t645[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t647 = FSM_dct_8x8_stage_2_0_t627;
    FSM_dct_8x8_stage_2_0_t647[FSM_dct_8x8_stage_2_0_t632 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t646;
    FSM_dct_8x8_stage_2_0_t648 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_2_0_t649 = FSM_dct_8x8_stage_2_0_t648[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t650 = FSM_dct_8x8_stage_2_0_t649 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_2_0_t651 = FSM_dct_8x8_stage_2_0_t650[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t652 = FSM_dct_8x8_stage_2_0_t651[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t653 = FSM_dct_8x8_stage_2_0_t647;
    FSM_dct_8x8_stage_2_0_t653[FSM_dct_8x8_stage_2_0_t652 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t638 - FSM_dct_8x8_stage_2_0_t644;
    FSM_dct_8x8_stage_2_0_t654 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_2_0_t655 = FSM_dct_8x8_stage_2_0_t654[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t656 = FSM_dct_8x8_stage_2_0_t655 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_2_0_t657 = FSM_dct_8x8_stage_2_0_t656[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t658 = FSM_dct_8x8_stage_2_0_t657[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t659 = FSM_dct_8x8_stage_2_0_t653;
    FSM_dct_8x8_stage_2_0_t659[FSM_dct_8x8_stage_2_0_t658 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t618 - FSM_dct_8x8_stage_2_0_t624;
    FSM_dct_8x8_stage_2_0_t660 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_2_0_t661 = FSM_dct_8x8_stage_2_0_t660[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t662 = FSM_dct_8x8_stage_2_0_t661 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_2_0_t663 = FSM_dct_8x8_stage_2_0_t662[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t664 = FSM_dct_8x8_stage_2_0_t663[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t665 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_2_0_t666 = FSM_dct_8x8_stage_2_0_t665[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t667 = FSM_dct_8x8_stage_2_0_t666 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_2_0_t668 = FSM_dct_8x8_stage_2_0_t667[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t669 = FSM_dct_8x8_stage_2_0_t668[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t670 = i_data_in[FSM_dct_8x8_stage_2_0_t669 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t671 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_2_0_t672 = FSM_dct_8x8_stage_2_0_t671[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t673 = FSM_dct_8x8_stage_2_0_t672 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_2_0_t674 = FSM_dct_8x8_stage_2_0_t673[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t675 = FSM_dct_8x8_stage_2_0_t674[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t676 = i_data_in[FSM_dct_8x8_stage_2_0_t675 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t677 = FSM_dct_8x8_stage_2_0_t670 + FSM_dct_8x8_stage_2_0_t676;
    FSM_dct_8x8_stage_2_0_t678 = FSM_dct_8x8_stage_2_0_t677[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t679 = FSM_dct_8x8_stage_2_0_t659;
    FSM_dct_8x8_stage_2_0_t679[FSM_dct_8x8_stage_2_0_t664 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t678;
    FSM_dct_8x8_stage_2_0_t680 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_2_0_t681 = FSM_dct_8x8_stage_2_0_t680[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t682 = FSM_dct_8x8_stage_2_0_t681 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_2_0_t683 = FSM_dct_8x8_stage_2_0_t682[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t684 = FSM_dct_8x8_stage_2_0_t683[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t685 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_2_0_t686 = FSM_dct_8x8_stage_2_0_t685[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t687 = FSM_dct_8x8_stage_2_0_t686 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_2_0_t688 = FSM_dct_8x8_stage_2_0_t687[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t689 = FSM_dct_8x8_stage_2_0_t688[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t690 = i_data_in[FSM_dct_8x8_stage_2_0_t689 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t691 = FSM_dct_8x8_stage_2_0_t676 + FSM_dct_8x8_stage_2_0_t690;
    FSM_dct_8x8_stage_2_0_t692 = FSM_dct_8x8_stage_2_0_t691[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t693 = FSM_dct_8x8_stage_2_0_t679;
    FSM_dct_8x8_stage_2_0_t693[FSM_dct_8x8_stage_2_0_t684 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t692;
    FSM_dct_8x8_stage_2_0_t694 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_2_0_t695 = FSM_dct_8x8_stage_2_0_t694[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t696 = FSM_dct_8x8_stage_2_0_t695 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_2_0_t697 = FSM_dct_8x8_stage_2_0_t696[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t698 = FSM_dct_8x8_stage_2_0_t697[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t699 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_2_0_t700 = FSM_dct_8x8_stage_2_0_t699[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t701 = FSM_dct_8x8_stage_2_0_t700 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_2_0_t702 = FSM_dct_8x8_stage_2_0_t701[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t703 = FSM_dct_8x8_stage_2_0_t702[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t704 = i_data_in[FSM_dct_8x8_stage_2_0_t703 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t705 = FSM_dct_8x8_stage_2_0_t690 + FSM_dct_8x8_stage_2_0_t704;
    FSM_dct_8x8_stage_2_0_t706 = FSM_dct_8x8_stage_2_0_t705[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t707 = FSM_dct_8x8_stage_2_0_t693;
    FSM_dct_8x8_stage_2_0_t707[FSM_dct_8x8_stage_2_0_t698 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t706;
    FSM_dct_8x8_stage_2_0_t708 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_2_0_t709 = FSM_dct_8x8_stage_2_0_t708[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t710 = FSM_dct_8x8_stage_2_0_t709 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_2_0_t711 = FSM_dct_8x8_stage_2_0_t710[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t712 = FSM_dct_8x8_stage_2_0_t711[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t713 = FSM_dct_8x8_stage_2_0_t707;
    FSM_dct_8x8_stage_2_0_t713[FSM_dct_8x8_stage_2_0_t712 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t704;
    FSM_dct_8x8_stage_2_0_t714 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_2_0_t715 = FSM_dct_8x8_stage_2_0_t714[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t716 = FSM_dct_8x8_stage_2_0_t715[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t717 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_2_0_t718 = FSM_dct_8x8_stage_2_0_t717[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t719 = FSM_dct_8x8_stage_2_0_t718[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t720 = i_data_in[FSM_dct_8x8_stage_2_0_t719 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t721 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_2_0_t722 = FSM_dct_8x8_stage_2_0_t721[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t723 = FSM_dct_8x8_stage_2_0_t722 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_2_0_t724 = FSM_dct_8x8_stage_2_0_t723[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t725 = FSM_dct_8x8_stage_2_0_t724[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t726 = i_data_in[FSM_dct_8x8_stage_2_0_t725 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t727 = FSM_dct_8x8_stage_2_0_t720 + FSM_dct_8x8_stage_2_0_t726;
    FSM_dct_8x8_stage_2_0_t728 = FSM_dct_8x8_stage_2_0_t727[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t729 = FSM_dct_8x8_stage_2_0_t713;
    FSM_dct_8x8_stage_2_0_t729[FSM_dct_8x8_stage_2_0_t716 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t728;
    FSM_dct_8x8_stage_2_0_t730 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_2_0_t731 = FSM_dct_8x8_stage_2_0_t730[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t732 = FSM_dct_8x8_stage_2_0_t731 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_2_0_t733 = FSM_dct_8x8_stage_2_0_t732[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t734 = FSM_dct_8x8_stage_2_0_t733[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t735 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_2_0_t736 = FSM_dct_8x8_stage_2_0_t735[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t737 = FSM_dct_8x8_stage_2_0_t736 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_2_0_t738 = FSM_dct_8x8_stage_2_0_t737[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t739 = FSM_dct_8x8_stage_2_0_t738[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t740 = i_data_in[FSM_dct_8x8_stage_2_0_t739 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t741 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_2_0_t742 = FSM_dct_8x8_stage_2_0_t741[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t743 = FSM_dct_8x8_stage_2_0_t742 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_2_0_t744 = FSM_dct_8x8_stage_2_0_t743[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t745 = FSM_dct_8x8_stage_2_0_t744[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t746 = i_data_in[FSM_dct_8x8_stage_2_0_t745 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t747 = FSM_dct_8x8_stage_2_0_t740 + FSM_dct_8x8_stage_2_0_t746;
    FSM_dct_8x8_stage_2_0_t748 = FSM_dct_8x8_stage_2_0_t747[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t749 = FSM_dct_8x8_stage_2_0_t729;
    FSM_dct_8x8_stage_2_0_t749[FSM_dct_8x8_stage_2_0_t734 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t748;
    FSM_dct_8x8_stage_2_0_t750 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_2_0_t751 = FSM_dct_8x8_stage_2_0_t750[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t752 = FSM_dct_8x8_stage_2_0_t751 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_2_0_t753 = FSM_dct_8x8_stage_2_0_t752[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t754 = FSM_dct_8x8_stage_2_0_t753[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t755 = FSM_dct_8x8_stage_2_0_t749;
    FSM_dct_8x8_stage_2_0_t755[FSM_dct_8x8_stage_2_0_t754 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t740 - FSM_dct_8x8_stage_2_0_t746;
    FSM_dct_8x8_stage_2_0_t756 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_2_0_t757 = FSM_dct_8x8_stage_2_0_t756[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t758 = FSM_dct_8x8_stage_2_0_t757 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_2_0_t759 = FSM_dct_8x8_stage_2_0_t758[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t760 = FSM_dct_8x8_stage_2_0_t759[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t761 = FSM_dct_8x8_stage_2_0_t755;
    FSM_dct_8x8_stage_2_0_t761[FSM_dct_8x8_stage_2_0_t760 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t720 - FSM_dct_8x8_stage_2_0_t726;
    FSM_dct_8x8_stage_2_0_t762 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_2_0_t763 = FSM_dct_8x8_stage_2_0_t762[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t764 = FSM_dct_8x8_stage_2_0_t763 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_2_0_t765 = FSM_dct_8x8_stage_2_0_t764[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t766 = FSM_dct_8x8_stage_2_0_t765[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t767 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_2_0_t768 = FSM_dct_8x8_stage_2_0_t767[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t769 = FSM_dct_8x8_stage_2_0_t768 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_2_0_t770 = FSM_dct_8x8_stage_2_0_t769[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t771 = FSM_dct_8x8_stage_2_0_t770[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t772 = i_data_in[FSM_dct_8x8_stage_2_0_t771 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t773 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_2_0_t774 = FSM_dct_8x8_stage_2_0_t773[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t775 = FSM_dct_8x8_stage_2_0_t774 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_2_0_t776 = FSM_dct_8x8_stage_2_0_t775[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t777 = FSM_dct_8x8_stage_2_0_t776[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t778 = i_data_in[FSM_dct_8x8_stage_2_0_t777 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t779 = FSM_dct_8x8_stage_2_0_t772 + FSM_dct_8x8_stage_2_0_t778;
    FSM_dct_8x8_stage_2_0_t780 = FSM_dct_8x8_stage_2_0_t779[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t781 = FSM_dct_8x8_stage_2_0_t761;
    FSM_dct_8x8_stage_2_0_t781[FSM_dct_8x8_stage_2_0_t766 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t780;
    FSM_dct_8x8_stage_2_0_t782 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_2_0_t783 = FSM_dct_8x8_stage_2_0_t782[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t784 = FSM_dct_8x8_stage_2_0_t783 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_2_0_t785 = FSM_dct_8x8_stage_2_0_t784[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t786 = FSM_dct_8x8_stage_2_0_t785[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t787 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_2_0_t788 = FSM_dct_8x8_stage_2_0_t787[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t789 = FSM_dct_8x8_stage_2_0_t788 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_2_0_t790 = FSM_dct_8x8_stage_2_0_t789[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t791 = FSM_dct_8x8_stage_2_0_t790[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t792 = i_data_in[FSM_dct_8x8_stage_2_0_t791 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t793 = FSM_dct_8x8_stage_2_0_t778 + FSM_dct_8x8_stage_2_0_t792;
    FSM_dct_8x8_stage_2_0_t794 = FSM_dct_8x8_stage_2_0_t793[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t795 = FSM_dct_8x8_stage_2_0_t781;
    FSM_dct_8x8_stage_2_0_t795[FSM_dct_8x8_stage_2_0_t786 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t794;
    FSM_dct_8x8_stage_2_0_t796 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_2_0_t797 = FSM_dct_8x8_stage_2_0_t796[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t798 = FSM_dct_8x8_stage_2_0_t797 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_2_0_t799 = FSM_dct_8x8_stage_2_0_t798[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t800 = FSM_dct_8x8_stage_2_0_t799[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t801 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_2_0_t802 = FSM_dct_8x8_stage_2_0_t801[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t803 = FSM_dct_8x8_stage_2_0_t802 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_2_0_t804 = FSM_dct_8x8_stage_2_0_t803[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t805 = FSM_dct_8x8_stage_2_0_t804[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t806 = i_data_in[FSM_dct_8x8_stage_2_0_t805 * 32 +: 32];
    FSM_dct_8x8_stage_2_0_t807 = FSM_dct_8x8_stage_2_0_t792 + FSM_dct_8x8_stage_2_0_t806;
    FSM_dct_8x8_stage_2_0_t808 = FSM_dct_8x8_stage_2_0_t807[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t809 = FSM_dct_8x8_stage_2_0_t795;
    FSM_dct_8x8_stage_2_0_t809[FSM_dct_8x8_stage_2_0_t800 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t808;
    FSM_dct_8x8_stage_2_0_t810 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_2_0_t811 = FSM_dct_8x8_stage_2_0_t810[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t812 = FSM_dct_8x8_stage_2_0_t811 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_2_0_t813 = FSM_dct_8x8_stage_2_0_t812[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_2_0_t814 = FSM_dct_8x8_stage_2_0_t813[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_2_0_t815 = FSM_dct_8x8_stage_2_0_t809;
    FSM_dct_8x8_stage_2_0_t815[FSM_dct_8x8_stage_2_0_t814 * 32 +: 32] = FSM_dct_8x8_stage_2_0_t806;
end

assign FSM_dct_8x8_stage_2_0_in_ready = 1'b1;

always @(posedge clk) begin
    FSM_dct_8x8_stage_2_0_st_dummy_reg <= FSM_dct_8x8_stage_2_0_st_dummy_reg;
    if (rst) begin
        FSM_dct_8x8_stage_2_0_st_dummy_reg <= 32'b0;
    end
end
/* End submodules of dct_8x8_stage_2 */
/* End module dct_8x8_stage_2 */
endgenerate
endmodule
