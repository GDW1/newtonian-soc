`timescale 1ns / 1ps

module dct_8x8_stage_1_inner
(
    input wire clk,
    input wire rst,
    input wire [2048-1:0] i_data_in,
    input wire i_valid,
    output wire i_ready,
    output wire [2048-1:0] o_data_out,
    output wire o_valid,
    input wire o_ready
);

generate
/*
    Begin module dct_8x8_stage_1
*/
/*
    Wires declared by dct_8x8_stage_1
*/
wire FSM_dct_8x8_stage_1_0_in_ready;
wire FSM_dct_8x8_stage_1_0_out_valid;
/* End wires declared by dct_8x8_stage_1 */

/*
    Submodules of dct_8x8_stage_1
*/
reg [32-1:0] FSM_dct_8x8_stage_1_0_st_dummy_reg = 32'b0;

reg [64-1:0] FSM_dct_8x8_stage_1_0_t0;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t1;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t2;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t3;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t4;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t5;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t6;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t7;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t8;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t9;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t10;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t11;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t12;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t13;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t14;
reg [2048-1:0] FSM_dct_8x8_stage_1_0_t15;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t16;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t17;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t18;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t19;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t20;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t21;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t22;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t23;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t24;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t25;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t26;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t27;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t28;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t29;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t30;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t31;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t32;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t33;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t34;
reg [2048-1:0] FSM_dct_8x8_stage_1_0_t35;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t36;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t37;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t38;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t39;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t40;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t41;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t42;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t43;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t44;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t45;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t46;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t47;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t48;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t49;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t50;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t51;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t52;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t53;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t54;
reg [2048-1:0] FSM_dct_8x8_stage_1_0_t55;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t56;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t57;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t58;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t59;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t60;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t61;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t62;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t63;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t64;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t65;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t66;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t67;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t68;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t69;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t70;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t71;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t72;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t73;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t74;
reg [2048-1:0] FSM_dct_8x8_stage_1_0_t75;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t76;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t77;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t78;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t79;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t80;
reg [2048-1:0] FSM_dct_8x8_stage_1_0_t81;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t82;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t83;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t84;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t85;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t86;
reg [2048-1:0] FSM_dct_8x8_stage_1_0_t87;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t88;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t89;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t90;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t91;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t92;
reg [2048-1:0] FSM_dct_8x8_stage_1_0_t93;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t94;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t95;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t96;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t97;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t98;
reg [2048-1:0] FSM_dct_8x8_stage_1_0_t99;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t100;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t101;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t102;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t103;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t104;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t105;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t106;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t107;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t108;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t109;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t110;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t111;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t112;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t113;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t114;
reg [2048-1:0] FSM_dct_8x8_stage_1_0_t115;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t116;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t117;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t118;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t119;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t120;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t121;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t122;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t123;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t124;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t125;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t126;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t127;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t128;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t129;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t130;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t131;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t132;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t133;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t134;
reg [2048-1:0] FSM_dct_8x8_stage_1_0_t135;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t136;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t137;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t138;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t139;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t140;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t141;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t142;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t143;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t144;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t145;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t146;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t147;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t148;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t149;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t150;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t151;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t152;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t153;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t154;
reg [2048-1:0] FSM_dct_8x8_stage_1_0_t155;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t156;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t157;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t158;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t159;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t160;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t161;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t162;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t163;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t164;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t165;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t166;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t167;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t168;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t169;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t170;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t171;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t172;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t173;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t174;
reg [2048-1:0] FSM_dct_8x8_stage_1_0_t175;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t176;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t177;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t178;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t179;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t180;
reg [2048-1:0] FSM_dct_8x8_stage_1_0_t181;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t182;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t183;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t184;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t185;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t186;
reg [2048-1:0] FSM_dct_8x8_stage_1_0_t187;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t188;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t189;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t190;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t191;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t192;
reg [2048-1:0] FSM_dct_8x8_stage_1_0_t193;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t194;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t195;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t196;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t197;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t198;
reg [2048-1:0] FSM_dct_8x8_stage_1_0_t199;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t200;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t201;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t202;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t203;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t204;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t205;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t206;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t207;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t208;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t209;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t210;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t211;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t212;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t213;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t214;
reg [2048-1:0] FSM_dct_8x8_stage_1_0_t215;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t216;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t217;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t218;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t219;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t220;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t221;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t222;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t223;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t224;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t225;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t226;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t227;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t228;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t229;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t230;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t231;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t232;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t233;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t234;
reg [2048-1:0] FSM_dct_8x8_stage_1_0_t235;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t236;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t237;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t238;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t239;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t240;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t241;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t242;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t243;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t244;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t245;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t246;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t247;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t248;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t249;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t250;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t251;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t252;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t253;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t254;
reg [2048-1:0] FSM_dct_8x8_stage_1_0_t255;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t256;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t257;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t258;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t259;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t260;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t261;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t262;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t263;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t264;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t265;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t266;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t267;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t268;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t269;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t270;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t271;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t272;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t273;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t274;
reg [2048-1:0] FSM_dct_8x8_stage_1_0_t275;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t276;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t277;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t278;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t279;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t280;
reg [2048-1:0] FSM_dct_8x8_stage_1_0_t281;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t282;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t283;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t284;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t285;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t286;
reg [2048-1:0] FSM_dct_8x8_stage_1_0_t287;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t288;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t289;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t290;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t291;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t292;
reg [2048-1:0] FSM_dct_8x8_stage_1_0_t293;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t294;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t295;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t296;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t297;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t298;
reg [2048-1:0] FSM_dct_8x8_stage_1_0_t299;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t300;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t301;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t302;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t303;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t304;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t305;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t306;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t307;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t308;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t309;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t310;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t311;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t312;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t313;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t314;
reg [2048-1:0] FSM_dct_8x8_stage_1_0_t315;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t316;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t317;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t318;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t319;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t320;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t321;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t322;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t323;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t324;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t325;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t326;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t327;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t328;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t329;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t330;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t331;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t332;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t333;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t334;
reg [2048-1:0] FSM_dct_8x8_stage_1_0_t335;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t336;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t337;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t338;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t339;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t340;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t341;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t342;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t343;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t344;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t345;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t346;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t347;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t348;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t349;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t350;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t351;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t352;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t353;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t354;
reg [2048-1:0] FSM_dct_8x8_stage_1_0_t355;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t356;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t357;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t358;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t359;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t360;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t361;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t362;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t363;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t364;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t365;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t366;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t367;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t368;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t369;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t370;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t371;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t372;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t373;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t374;
reg [2048-1:0] FSM_dct_8x8_stage_1_0_t375;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t376;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t377;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t378;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t379;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t380;
reg [2048-1:0] FSM_dct_8x8_stage_1_0_t381;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t382;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t383;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t384;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t385;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t386;
reg [2048-1:0] FSM_dct_8x8_stage_1_0_t387;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t388;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t389;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t390;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t391;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t392;
reg [2048-1:0] FSM_dct_8x8_stage_1_0_t393;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t394;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t395;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t396;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t397;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t398;
reg [2048-1:0] FSM_dct_8x8_stage_1_0_t399;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t400;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t401;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t402;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t403;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t404;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t405;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t406;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t407;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t408;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t409;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t410;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t411;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t412;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t413;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t414;
reg [2048-1:0] FSM_dct_8x8_stage_1_0_t415;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t416;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t417;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t418;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t419;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t420;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t421;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t422;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t423;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t424;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t425;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t426;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t427;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t428;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t429;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t430;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t431;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t432;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t433;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t434;
reg [2048-1:0] FSM_dct_8x8_stage_1_0_t435;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t436;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t437;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t438;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t439;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t440;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t441;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t442;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t443;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t444;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t445;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t446;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t447;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t448;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t449;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t450;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t451;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t452;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t453;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t454;
reg [2048-1:0] FSM_dct_8x8_stage_1_0_t455;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t456;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t457;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t458;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t459;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t460;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t461;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t462;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t463;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t464;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t465;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t466;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t467;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t468;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t469;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t470;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t471;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t472;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t473;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t474;
reg [2048-1:0] FSM_dct_8x8_stage_1_0_t475;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t476;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t477;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t478;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t479;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t480;
reg [2048-1:0] FSM_dct_8x8_stage_1_0_t481;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t482;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t483;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t484;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t485;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t486;
reg [2048-1:0] FSM_dct_8x8_stage_1_0_t487;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t488;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t489;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t490;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t491;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t492;
reg [2048-1:0] FSM_dct_8x8_stage_1_0_t493;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t494;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t495;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t496;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t497;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t498;
reg [2048-1:0] FSM_dct_8x8_stage_1_0_t499;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t500;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t501;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t502;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t503;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t504;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t505;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t506;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t507;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t508;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t509;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t510;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t511;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t512;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t513;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t514;
reg [2048-1:0] FSM_dct_8x8_stage_1_0_t515;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t516;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t517;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t518;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t519;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t520;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t521;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t522;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t523;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t524;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t525;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t526;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t527;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t528;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t529;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t530;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t531;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t532;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t533;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t534;
reg [2048-1:0] FSM_dct_8x8_stage_1_0_t535;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t536;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t537;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t538;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t539;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t540;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t541;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t542;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t543;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t544;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t545;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t546;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t547;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t548;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t549;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t550;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t551;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t552;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t553;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t554;
reg [2048-1:0] FSM_dct_8x8_stage_1_0_t555;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t556;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t557;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t558;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t559;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t560;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t561;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t562;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t563;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t564;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t565;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t566;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t567;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t568;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t569;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t570;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t571;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t572;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t573;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t574;
reg [2048-1:0] FSM_dct_8x8_stage_1_0_t575;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t576;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t577;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t578;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t579;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t580;
reg [2048-1:0] FSM_dct_8x8_stage_1_0_t581;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t582;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t583;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t584;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t585;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t586;
reg [2048-1:0] FSM_dct_8x8_stage_1_0_t587;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t588;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t589;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t590;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t591;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t592;
reg [2048-1:0] FSM_dct_8x8_stage_1_0_t593;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t594;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t595;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t596;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t597;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t598;
reg [2048-1:0] FSM_dct_8x8_stage_1_0_t599;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t600;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t601;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t602;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t603;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t604;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t605;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t606;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t607;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t608;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t609;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t610;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t611;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t612;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t613;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t614;
reg [2048-1:0] FSM_dct_8x8_stage_1_0_t615;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t616;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t617;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t618;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t619;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t620;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t621;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t622;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t623;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t624;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t625;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t626;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t627;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t628;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t629;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t630;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t631;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t632;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t633;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t634;
reg [2048-1:0] FSM_dct_8x8_stage_1_0_t635;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t636;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t637;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t638;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t639;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t640;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t641;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t642;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t643;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t644;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t645;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t646;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t647;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t648;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t649;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t650;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t651;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t652;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t653;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t654;
reg [2048-1:0] FSM_dct_8x8_stage_1_0_t655;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t656;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t657;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t658;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t659;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t660;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t661;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t662;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t663;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t664;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t665;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t666;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t667;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t668;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t669;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t670;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t671;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t672;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t673;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t674;
reg [2048-1:0] FSM_dct_8x8_stage_1_0_t675;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t676;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t677;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t678;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t679;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t680;
reg [2048-1:0] FSM_dct_8x8_stage_1_0_t681;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t682;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t683;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t684;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t685;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t686;
reg [2048-1:0] FSM_dct_8x8_stage_1_0_t687;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t688;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t689;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t690;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t691;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t692;
reg [2048-1:0] FSM_dct_8x8_stage_1_0_t693;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t694;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t695;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t696;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t697;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t698;
reg [2048-1:0] FSM_dct_8x8_stage_1_0_t699;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t700;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t701;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t702;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t703;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t704;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t705;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t706;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t707;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t708;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t709;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t710;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t711;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t712;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t713;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t714;
reg [2048-1:0] FSM_dct_8x8_stage_1_0_t715;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t716;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t717;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t718;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t719;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t720;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t721;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t722;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t723;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t724;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t725;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t726;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t727;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t728;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t729;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t730;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t731;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t732;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t733;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t734;
reg [2048-1:0] FSM_dct_8x8_stage_1_0_t735;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t736;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t737;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t738;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t739;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t740;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t741;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t742;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t743;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t744;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t745;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t746;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t747;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t748;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t749;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t750;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t751;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t752;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t753;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t754;
reg [2048-1:0] FSM_dct_8x8_stage_1_0_t755;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t756;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t757;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t758;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t759;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t760;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t761;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t762;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t763;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t764;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t765;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t766;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t767;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t768;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t769;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t770;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t771;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t772;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t773;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t774;
reg [2048-1:0] FSM_dct_8x8_stage_1_0_t775;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t776;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t777;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t778;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t779;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t780;
reg [2048-1:0] FSM_dct_8x8_stage_1_0_t781;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t782;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t783;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t784;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t785;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t786;
reg [2048-1:0] FSM_dct_8x8_stage_1_0_t787;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t788;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t789;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t790;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t791;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t792;
reg [2048-1:0] FSM_dct_8x8_stage_1_0_t793;
reg [64-1:0] FSM_dct_8x8_stage_1_0_t794;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t795;
reg [33-1:0] FSM_dct_8x8_stage_1_0_t796;
reg [32-1:0] FSM_dct_8x8_stage_1_0_t797;
reg [6-1:0] FSM_dct_8x8_stage_1_0_t798;
reg [2048-1:0] FSM_dct_8x8_stage_1_0_t799;

/*
    Wiring by dct_8x8_stage_1
*/
assign i_ready = FSM_dct_8x8_stage_1_0_in_ready;
assign o_data_out = FSM_dct_8x8_stage_1_0_t799;
assign o_valid = FSM_dct_8x8_stage_1_0_out_valid;
/* End wiring by dct_8x8_stage_1 */

assign FSM_dct_8x8_stage_1_0_out_valid = 1'b1;

initial begin
    FSM_dct_8x8_stage_1_0_t0 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_1_0_t1 = FSM_dct_8x8_stage_1_0_t0[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t2 = FSM_dct_8x8_stage_1_0_t1[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t3 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_1_0_t4 = FSM_dct_8x8_stage_1_0_t3[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t5 = FSM_dct_8x8_stage_1_0_t4[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t6 = i_data_in[FSM_dct_8x8_stage_1_0_t5 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t7 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_1_0_t8 = FSM_dct_8x8_stage_1_0_t7[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t9 = FSM_dct_8x8_stage_1_0_t8 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_1_0_t10 = FSM_dct_8x8_stage_1_0_t9[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t11 = FSM_dct_8x8_stage_1_0_t10[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t12 = i_data_in[FSM_dct_8x8_stage_1_0_t11 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t13 = FSM_dct_8x8_stage_1_0_t6 + FSM_dct_8x8_stage_1_0_t12;
    FSM_dct_8x8_stage_1_0_t14 = FSM_dct_8x8_stage_1_0_t13[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t15 = 2048'b0;
    FSM_dct_8x8_stage_1_0_t15[FSM_dct_8x8_stage_1_0_t2 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t14;
    FSM_dct_8x8_stage_1_0_t16 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_1_0_t17 = FSM_dct_8x8_stage_1_0_t16[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t18 = FSM_dct_8x8_stage_1_0_t17 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_1_0_t19 = FSM_dct_8x8_stage_1_0_t18[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t20 = FSM_dct_8x8_stage_1_0_t19[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t21 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_1_0_t22 = FSM_dct_8x8_stage_1_0_t21[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t23 = FSM_dct_8x8_stage_1_0_t22 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_1_0_t24 = FSM_dct_8x8_stage_1_0_t23[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t25 = FSM_dct_8x8_stage_1_0_t24[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t26 = i_data_in[FSM_dct_8x8_stage_1_0_t25 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t27 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_1_0_t28 = FSM_dct_8x8_stage_1_0_t27[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t29 = FSM_dct_8x8_stage_1_0_t28 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_1_0_t30 = FSM_dct_8x8_stage_1_0_t29[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t31 = FSM_dct_8x8_stage_1_0_t30[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t32 = i_data_in[FSM_dct_8x8_stage_1_0_t31 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t33 = FSM_dct_8x8_stage_1_0_t26 + FSM_dct_8x8_stage_1_0_t32;
    FSM_dct_8x8_stage_1_0_t34 = FSM_dct_8x8_stage_1_0_t33[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t35 = FSM_dct_8x8_stage_1_0_t15;
    FSM_dct_8x8_stage_1_0_t35[FSM_dct_8x8_stage_1_0_t20 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t34;
    FSM_dct_8x8_stage_1_0_t36 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_1_0_t37 = FSM_dct_8x8_stage_1_0_t36[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t38 = FSM_dct_8x8_stage_1_0_t37 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_1_0_t39 = FSM_dct_8x8_stage_1_0_t38[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t40 = FSM_dct_8x8_stage_1_0_t39[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t41 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_1_0_t42 = FSM_dct_8x8_stage_1_0_t41[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t43 = FSM_dct_8x8_stage_1_0_t42 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_1_0_t44 = FSM_dct_8x8_stage_1_0_t43[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t45 = FSM_dct_8x8_stage_1_0_t44[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t46 = i_data_in[FSM_dct_8x8_stage_1_0_t45 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t47 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_1_0_t48 = FSM_dct_8x8_stage_1_0_t47[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t49 = FSM_dct_8x8_stage_1_0_t48 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_1_0_t50 = FSM_dct_8x8_stage_1_0_t49[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t51 = FSM_dct_8x8_stage_1_0_t50[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t52 = i_data_in[FSM_dct_8x8_stage_1_0_t51 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t53 = FSM_dct_8x8_stage_1_0_t46 + FSM_dct_8x8_stage_1_0_t52;
    FSM_dct_8x8_stage_1_0_t54 = FSM_dct_8x8_stage_1_0_t53[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t55 = FSM_dct_8x8_stage_1_0_t35;
    FSM_dct_8x8_stage_1_0_t55[FSM_dct_8x8_stage_1_0_t40 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t54;
    FSM_dct_8x8_stage_1_0_t56 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_1_0_t57 = FSM_dct_8x8_stage_1_0_t56[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t58 = FSM_dct_8x8_stage_1_0_t57 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_1_0_t59 = FSM_dct_8x8_stage_1_0_t58[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t60 = FSM_dct_8x8_stage_1_0_t59[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t61 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_1_0_t62 = FSM_dct_8x8_stage_1_0_t61[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t63 = FSM_dct_8x8_stage_1_0_t62 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_1_0_t64 = FSM_dct_8x8_stage_1_0_t63[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t65 = FSM_dct_8x8_stage_1_0_t64[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t66 = i_data_in[FSM_dct_8x8_stage_1_0_t65 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t67 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_1_0_t68 = FSM_dct_8x8_stage_1_0_t67[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t69 = FSM_dct_8x8_stage_1_0_t68 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_1_0_t70 = FSM_dct_8x8_stage_1_0_t69[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t71 = FSM_dct_8x8_stage_1_0_t70[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t72 = i_data_in[FSM_dct_8x8_stage_1_0_t71 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t73 = FSM_dct_8x8_stage_1_0_t66 + FSM_dct_8x8_stage_1_0_t72;
    FSM_dct_8x8_stage_1_0_t74 = FSM_dct_8x8_stage_1_0_t73[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t75 = FSM_dct_8x8_stage_1_0_t55;
    FSM_dct_8x8_stage_1_0_t75[FSM_dct_8x8_stage_1_0_t60 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t74;
    FSM_dct_8x8_stage_1_0_t76 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_1_0_t77 = FSM_dct_8x8_stage_1_0_t76[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t78 = FSM_dct_8x8_stage_1_0_t77 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_1_0_t79 = FSM_dct_8x8_stage_1_0_t78[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t80 = FSM_dct_8x8_stage_1_0_t79[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t81 = FSM_dct_8x8_stage_1_0_t75;
    FSM_dct_8x8_stage_1_0_t81[FSM_dct_8x8_stage_1_0_t80 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t66 - FSM_dct_8x8_stage_1_0_t72;
    FSM_dct_8x8_stage_1_0_t82 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_1_0_t83 = FSM_dct_8x8_stage_1_0_t82[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t84 = FSM_dct_8x8_stage_1_0_t83 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_1_0_t85 = FSM_dct_8x8_stage_1_0_t84[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t86 = FSM_dct_8x8_stage_1_0_t85[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t87 = FSM_dct_8x8_stage_1_0_t81;
    FSM_dct_8x8_stage_1_0_t87[FSM_dct_8x8_stage_1_0_t86 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t46 - FSM_dct_8x8_stage_1_0_t52;
    FSM_dct_8x8_stage_1_0_t88 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_1_0_t89 = FSM_dct_8x8_stage_1_0_t88[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t90 = FSM_dct_8x8_stage_1_0_t89 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_1_0_t91 = FSM_dct_8x8_stage_1_0_t90[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t92 = FSM_dct_8x8_stage_1_0_t91[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t93 = FSM_dct_8x8_stage_1_0_t87;
    FSM_dct_8x8_stage_1_0_t93[FSM_dct_8x8_stage_1_0_t92 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t26 - FSM_dct_8x8_stage_1_0_t32;
    FSM_dct_8x8_stage_1_0_t94 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_1_0_t95 = FSM_dct_8x8_stage_1_0_t94[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t96 = FSM_dct_8x8_stage_1_0_t95 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_1_0_t97 = FSM_dct_8x8_stage_1_0_t96[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t98 = FSM_dct_8x8_stage_1_0_t97[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t99 = FSM_dct_8x8_stage_1_0_t93;
    FSM_dct_8x8_stage_1_0_t99[FSM_dct_8x8_stage_1_0_t98 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t6 - FSM_dct_8x8_stage_1_0_t12;
    FSM_dct_8x8_stage_1_0_t100 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_1_0_t101 = FSM_dct_8x8_stage_1_0_t100[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t102 = FSM_dct_8x8_stage_1_0_t101[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t103 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_1_0_t104 = FSM_dct_8x8_stage_1_0_t103[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t105 = FSM_dct_8x8_stage_1_0_t104[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t106 = i_data_in[FSM_dct_8x8_stage_1_0_t105 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t107 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_1_0_t108 = FSM_dct_8x8_stage_1_0_t107[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t109 = FSM_dct_8x8_stage_1_0_t108 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_1_0_t110 = FSM_dct_8x8_stage_1_0_t109[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t111 = FSM_dct_8x8_stage_1_0_t110[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t112 = i_data_in[FSM_dct_8x8_stage_1_0_t111 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t113 = FSM_dct_8x8_stage_1_0_t106 + FSM_dct_8x8_stage_1_0_t112;
    FSM_dct_8x8_stage_1_0_t114 = FSM_dct_8x8_stage_1_0_t113[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t115 = FSM_dct_8x8_stage_1_0_t99;
    FSM_dct_8x8_stage_1_0_t115[FSM_dct_8x8_stage_1_0_t102 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t114;
    FSM_dct_8x8_stage_1_0_t116 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_1_0_t117 = FSM_dct_8x8_stage_1_0_t116[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t118 = FSM_dct_8x8_stage_1_0_t117 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_1_0_t119 = FSM_dct_8x8_stage_1_0_t118[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t120 = FSM_dct_8x8_stage_1_0_t119[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t121 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_1_0_t122 = FSM_dct_8x8_stage_1_0_t121[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t123 = FSM_dct_8x8_stage_1_0_t122 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_1_0_t124 = FSM_dct_8x8_stage_1_0_t123[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t125 = FSM_dct_8x8_stage_1_0_t124[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t126 = i_data_in[FSM_dct_8x8_stage_1_0_t125 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t127 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_1_0_t128 = FSM_dct_8x8_stage_1_0_t127[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t129 = FSM_dct_8x8_stage_1_0_t128 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_1_0_t130 = FSM_dct_8x8_stage_1_0_t129[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t131 = FSM_dct_8x8_stage_1_0_t130[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t132 = i_data_in[FSM_dct_8x8_stage_1_0_t131 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t133 = FSM_dct_8x8_stage_1_0_t126 + FSM_dct_8x8_stage_1_0_t132;
    FSM_dct_8x8_stage_1_0_t134 = FSM_dct_8x8_stage_1_0_t133[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t135 = FSM_dct_8x8_stage_1_0_t115;
    FSM_dct_8x8_stage_1_0_t135[FSM_dct_8x8_stage_1_0_t120 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t134;
    FSM_dct_8x8_stage_1_0_t136 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_1_0_t137 = FSM_dct_8x8_stage_1_0_t136[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t138 = FSM_dct_8x8_stage_1_0_t137 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_1_0_t139 = FSM_dct_8x8_stage_1_0_t138[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t140 = FSM_dct_8x8_stage_1_0_t139[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t141 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_1_0_t142 = FSM_dct_8x8_stage_1_0_t141[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t143 = FSM_dct_8x8_stage_1_0_t142 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_1_0_t144 = FSM_dct_8x8_stage_1_0_t143[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t145 = FSM_dct_8x8_stage_1_0_t144[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t146 = i_data_in[FSM_dct_8x8_stage_1_0_t145 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t147 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_1_0_t148 = FSM_dct_8x8_stage_1_0_t147[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t149 = FSM_dct_8x8_stage_1_0_t148 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_1_0_t150 = FSM_dct_8x8_stage_1_0_t149[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t151 = FSM_dct_8x8_stage_1_0_t150[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t152 = i_data_in[FSM_dct_8x8_stage_1_0_t151 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t153 = FSM_dct_8x8_stage_1_0_t146 + FSM_dct_8x8_stage_1_0_t152;
    FSM_dct_8x8_stage_1_0_t154 = FSM_dct_8x8_stage_1_0_t153[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t155 = FSM_dct_8x8_stage_1_0_t135;
    FSM_dct_8x8_stage_1_0_t155[FSM_dct_8x8_stage_1_0_t140 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t154;
    FSM_dct_8x8_stage_1_0_t156 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_1_0_t157 = FSM_dct_8x8_stage_1_0_t156[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t158 = FSM_dct_8x8_stage_1_0_t157 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_1_0_t159 = FSM_dct_8x8_stage_1_0_t158[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t160 = FSM_dct_8x8_stage_1_0_t159[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t161 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_1_0_t162 = FSM_dct_8x8_stage_1_0_t161[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t163 = FSM_dct_8x8_stage_1_0_t162 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_1_0_t164 = FSM_dct_8x8_stage_1_0_t163[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t165 = FSM_dct_8x8_stage_1_0_t164[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t166 = i_data_in[FSM_dct_8x8_stage_1_0_t165 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t167 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_1_0_t168 = FSM_dct_8x8_stage_1_0_t167[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t169 = FSM_dct_8x8_stage_1_0_t168 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_1_0_t170 = FSM_dct_8x8_stage_1_0_t169[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t171 = FSM_dct_8x8_stage_1_0_t170[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t172 = i_data_in[FSM_dct_8x8_stage_1_0_t171 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t173 = FSM_dct_8x8_stage_1_0_t166 + FSM_dct_8x8_stage_1_0_t172;
    FSM_dct_8x8_stage_1_0_t174 = FSM_dct_8x8_stage_1_0_t173[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t175 = FSM_dct_8x8_stage_1_0_t155;
    FSM_dct_8x8_stage_1_0_t175[FSM_dct_8x8_stage_1_0_t160 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t174;
    FSM_dct_8x8_stage_1_0_t176 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_1_0_t177 = FSM_dct_8x8_stage_1_0_t176[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t178 = FSM_dct_8x8_stage_1_0_t177 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_1_0_t179 = FSM_dct_8x8_stage_1_0_t178[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t180 = FSM_dct_8x8_stage_1_0_t179[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t181 = FSM_dct_8x8_stage_1_0_t175;
    FSM_dct_8x8_stage_1_0_t181[FSM_dct_8x8_stage_1_0_t180 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t166 - FSM_dct_8x8_stage_1_0_t172;
    FSM_dct_8x8_stage_1_0_t182 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_1_0_t183 = FSM_dct_8x8_stage_1_0_t182[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t184 = FSM_dct_8x8_stage_1_0_t183 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_1_0_t185 = FSM_dct_8x8_stage_1_0_t184[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t186 = FSM_dct_8x8_stage_1_0_t185[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t187 = FSM_dct_8x8_stage_1_0_t181;
    FSM_dct_8x8_stage_1_0_t187[FSM_dct_8x8_stage_1_0_t186 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t146 - FSM_dct_8x8_stage_1_0_t152;
    FSM_dct_8x8_stage_1_0_t188 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_1_0_t189 = FSM_dct_8x8_stage_1_0_t188[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t190 = FSM_dct_8x8_stage_1_0_t189 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_1_0_t191 = FSM_dct_8x8_stage_1_0_t190[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t192 = FSM_dct_8x8_stage_1_0_t191[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t193 = FSM_dct_8x8_stage_1_0_t187;
    FSM_dct_8x8_stage_1_0_t193[FSM_dct_8x8_stage_1_0_t192 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t126 - FSM_dct_8x8_stage_1_0_t132;
    FSM_dct_8x8_stage_1_0_t194 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_1_0_t195 = FSM_dct_8x8_stage_1_0_t194[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t196 = FSM_dct_8x8_stage_1_0_t195 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_1_0_t197 = FSM_dct_8x8_stage_1_0_t196[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t198 = FSM_dct_8x8_stage_1_0_t197[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t199 = FSM_dct_8x8_stage_1_0_t193;
    FSM_dct_8x8_stage_1_0_t199[FSM_dct_8x8_stage_1_0_t198 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t106 - FSM_dct_8x8_stage_1_0_t112;
    FSM_dct_8x8_stage_1_0_t200 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_1_0_t201 = FSM_dct_8x8_stage_1_0_t200[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t202 = FSM_dct_8x8_stage_1_0_t201[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t203 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_1_0_t204 = FSM_dct_8x8_stage_1_0_t203[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t205 = FSM_dct_8x8_stage_1_0_t204[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t206 = i_data_in[FSM_dct_8x8_stage_1_0_t205 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t207 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_1_0_t208 = FSM_dct_8x8_stage_1_0_t207[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t209 = FSM_dct_8x8_stage_1_0_t208 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_1_0_t210 = FSM_dct_8x8_stage_1_0_t209[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t211 = FSM_dct_8x8_stage_1_0_t210[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t212 = i_data_in[FSM_dct_8x8_stage_1_0_t211 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t213 = FSM_dct_8x8_stage_1_0_t206 + FSM_dct_8x8_stage_1_0_t212;
    FSM_dct_8x8_stage_1_0_t214 = FSM_dct_8x8_stage_1_0_t213[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t215 = FSM_dct_8x8_stage_1_0_t199;
    FSM_dct_8x8_stage_1_0_t215[FSM_dct_8x8_stage_1_0_t202 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t214;
    FSM_dct_8x8_stage_1_0_t216 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_1_0_t217 = FSM_dct_8x8_stage_1_0_t216[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t218 = FSM_dct_8x8_stage_1_0_t217 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_1_0_t219 = FSM_dct_8x8_stage_1_0_t218[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t220 = FSM_dct_8x8_stage_1_0_t219[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t221 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_1_0_t222 = FSM_dct_8x8_stage_1_0_t221[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t223 = FSM_dct_8x8_stage_1_0_t222 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_1_0_t224 = FSM_dct_8x8_stage_1_0_t223[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t225 = FSM_dct_8x8_stage_1_0_t224[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t226 = i_data_in[FSM_dct_8x8_stage_1_0_t225 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t227 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_1_0_t228 = FSM_dct_8x8_stage_1_0_t227[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t229 = FSM_dct_8x8_stage_1_0_t228 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_1_0_t230 = FSM_dct_8x8_stage_1_0_t229[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t231 = FSM_dct_8x8_stage_1_0_t230[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t232 = i_data_in[FSM_dct_8x8_stage_1_0_t231 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t233 = FSM_dct_8x8_stage_1_0_t226 + FSM_dct_8x8_stage_1_0_t232;
    FSM_dct_8x8_stage_1_0_t234 = FSM_dct_8x8_stage_1_0_t233[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t235 = FSM_dct_8x8_stage_1_0_t215;
    FSM_dct_8x8_stage_1_0_t235[FSM_dct_8x8_stage_1_0_t220 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t234;
    FSM_dct_8x8_stage_1_0_t236 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_1_0_t237 = FSM_dct_8x8_stage_1_0_t236[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t238 = FSM_dct_8x8_stage_1_0_t237 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_1_0_t239 = FSM_dct_8x8_stage_1_0_t238[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t240 = FSM_dct_8x8_stage_1_0_t239[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t241 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_1_0_t242 = FSM_dct_8x8_stage_1_0_t241[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t243 = FSM_dct_8x8_stage_1_0_t242 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_1_0_t244 = FSM_dct_8x8_stage_1_0_t243[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t245 = FSM_dct_8x8_stage_1_0_t244[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t246 = i_data_in[FSM_dct_8x8_stage_1_0_t245 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t247 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_1_0_t248 = FSM_dct_8x8_stage_1_0_t247[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t249 = FSM_dct_8x8_stage_1_0_t248 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_1_0_t250 = FSM_dct_8x8_stage_1_0_t249[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t251 = FSM_dct_8x8_stage_1_0_t250[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t252 = i_data_in[FSM_dct_8x8_stage_1_0_t251 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t253 = FSM_dct_8x8_stage_1_0_t246 + FSM_dct_8x8_stage_1_0_t252;
    FSM_dct_8x8_stage_1_0_t254 = FSM_dct_8x8_stage_1_0_t253[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t255 = FSM_dct_8x8_stage_1_0_t235;
    FSM_dct_8x8_stage_1_0_t255[FSM_dct_8x8_stage_1_0_t240 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t254;
    FSM_dct_8x8_stage_1_0_t256 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_1_0_t257 = FSM_dct_8x8_stage_1_0_t256[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t258 = FSM_dct_8x8_stage_1_0_t257 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_1_0_t259 = FSM_dct_8x8_stage_1_0_t258[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t260 = FSM_dct_8x8_stage_1_0_t259[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t261 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_1_0_t262 = FSM_dct_8x8_stage_1_0_t261[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t263 = FSM_dct_8x8_stage_1_0_t262 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_1_0_t264 = FSM_dct_8x8_stage_1_0_t263[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t265 = FSM_dct_8x8_stage_1_0_t264[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t266 = i_data_in[FSM_dct_8x8_stage_1_0_t265 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t267 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_1_0_t268 = FSM_dct_8x8_stage_1_0_t267[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t269 = FSM_dct_8x8_stage_1_0_t268 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_1_0_t270 = FSM_dct_8x8_stage_1_0_t269[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t271 = FSM_dct_8x8_stage_1_0_t270[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t272 = i_data_in[FSM_dct_8x8_stage_1_0_t271 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t273 = FSM_dct_8x8_stage_1_0_t266 + FSM_dct_8x8_stage_1_0_t272;
    FSM_dct_8x8_stage_1_0_t274 = FSM_dct_8x8_stage_1_0_t273[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t275 = FSM_dct_8x8_stage_1_0_t255;
    FSM_dct_8x8_stage_1_0_t275[FSM_dct_8x8_stage_1_0_t260 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t274;
    FSM_dct_8x8_stage_1_0_t276 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_1_0_t277 = FSM_dct_8x8_stage_1_0_t276[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t278 = FSM_dct_8x8_stage_1_0_t277 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_1_0_t279 = FSM_dct_8x8_stage_1_0_t278[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t280 = FSM_dct_8x8_stage_1_0_t279[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t281 = FSM_dct_8x8_stage_1_0_t275;
    FSM_dct_8x8_stage_1_0_t281[FSM_dct_8x8_stage_1_0_t280 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t266 - FSM_dct_8x8_stage_1_0_t272;
    FSM_dct_8x8_stage_1_0_t282 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_1_0_t283 = FSM_dct_8x8_stage_1_0_t282[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t284 = FSM_dct_8x8_stage_1_0_t283 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_1_0_t285 = FSM_dct_8x8_stage_1_0_t284[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t286 = FSM_dct_8x8_stage_1_0_t285[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t287 = FSM_dct_8x8_stage_1_0_t281;
    FSM_dct_8x8_stage_1_0_t287[FSM_dct_8x8_stage_1_0_t286 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t246 - FSM_dct_8x8_stage_1_0_t252;
    FSM_dct_8x8_stage_1_0_t288 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_1_0_t289 = FSM_dct_8x8_stage_1_0_t288[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t290 = FSM_dct_8x8_stage_1_0_t289 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_1_0_t291 = FSM_dct_8x8_stage_1_0_t290[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t292 = FSM_dct_8x8_stage_1_0_t291[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t293 = FSM_dct_8x8_stage_1_0_t287;
    FSM_dct_8x8_stage_1_0_t293[FSM_dct_8x8_stage_1_0_t292 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t226 - FSM_dct_8x8_stage_1_0_t232;
    FSM_dct_8x8_stage_1_0_t294 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_1_0_t295 = FSM_dct_8x8_stage_1_0_t294[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t296 = FSM_dct_8x8_stage_1_0_t295 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_1_0_t297 = FSM_dct_8x8_stage_1_0_t296[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t298 = FSM_dct_8x8_stage_1_0_t297[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t299 = FSM_dct_8x8_stage_1_0_t293;
    FSM_dct_8x8_stage_1_0_t299[FSM_dct_8x8_stage_1_0_t298 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t206 - FSM_dct_8x8_stage_1_0_t212;
    FSM_dct_8x8_stage_1_0_t300 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_1_0_t301 = FSM_dct_8x8_stage_1_0_t300[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t302 = FSM_dct_8x8_stage_1_0_t301[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t303 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_1_0_t304 = FSM_dct_8x8_stage_1_0_t303[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t305 = FSM_dct_8x8_stage_1_0_t304[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t306 = i_data_in[FSM_dct_8x8_stage_1_0_t305 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t307 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_1_0_t308 = FSM_dct_8x8_stage_1_0_t307[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t309 = FSM_dct_8x8_stage_1_0_t308 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_1_0_t310 = FSM_dct_8x8_stage_1_0_t309[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t311 = FSM_dct_8x8_stage_1_0_t310[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t312 = i_data_in[FSM_dct_8x8_stage_1_0_t311 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t313 = FSM_dct_8x8_stage_1_0_t306 + FSM_dct_8x8_stage_1_0_t312;
    FSM_dct_8x8_stage_1_0_t314 = FSM_dct_8x8_stage_1_0_t313[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t315 = FSM_dct_8x8_stage_1_0_t299;
    FSM_dct_8x8_stage_1_0_t315[FSM_dct_8x8_stage_1_0_t302 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t314;
    FSM_dct_8x8_stage_1_0_t316 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_1_0_t317 = FSM_dct_8x8_stage_1_0_t316[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t318 = FSM_dct_8x8_stage_1_0_t317 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_1_0_t319 = FSM_dct_8x8_stage_1_0_t318[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t320 = FSM_dct_8x8_stage_1_0_t319[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t321 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_1_0_t322 = FSM_dct_8x8_stage_1_0_t321[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t323 = FSM_dct_8x8_stage_1_0_t322 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_1_0_t324 = FSM_dct_8x8_stage_1_0_t323[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t325 = FSM_dct_8x8_stage_1_0_t324[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t326 = i_data_in[FSM_dct_8x8_stage_1_0_t325 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t327 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_1_0_t328 = FSM_dct_8x8_stage_1_0_t327[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t329 = FSM_dct_8x8_stage_1_0_t328 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_1_0_t330 = FSM_dct_8x8_stage_1_0_t329[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t331 = FSM_dct_8x8_stage_1_0_t330[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t332 = i_data_in[FSM_dct_8x8_stage_1_0_t331 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t333 = FSM_dct_8x8_stage_1_0_t326 + FSM_dct_8x8_stage_1_0_t332;
    FSM_dct_8x8_stage_1_0_t334 = FSM_dct_8x8_stage_1_0_t333[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t335 = FSM_dct_8x8_stage_1_0_t315;
    FSM_dct_8x8_stage_1_0_t335[FSM_dct_8x8_stage_1_0_t320 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t334;
    FSM_dct_8x8_stage_1_0_t336 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_1_0_t337 = FSM_dct_8x8_stage_1_0_t336[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t338 = FSM_dct_8x8_stage_1_0_t337 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_1_0_t339 = FSM_dct_8x8_stage_1_0_t338[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t340 = FSM_dct_8x8_stage_1_0_t339[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t341 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_1_0_t342 = FSM_dct_8x8_stage_1_0_t341[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t343 = FSM_dct_8x8_stage_1_0_t342 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_1_0_t344 = FSM_dct_8x8_stage_1_0_t343[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t345 = FSM_dct_8x8_stage_1_0_t344[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t346 = i_data_in[FSM_dct_8x8_stage_1_0_t345 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t347 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_1_0_t348 = FSM_dct_8x8_stage_1_0_t347[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t349 = FSM_dct_8x8_stage_1_0_t348 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_1_0_t350 = FSM_dct_8x8_stage_1_0_t349[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t351 = FSM_dct_8x8_stage_1_0_t350[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t352 = i_data_in[FSM_dct_8x8_stage_1_0_t351 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t353 = FSM_dct_8x8_stage_1_0_t346 + FSM_dct_8x8_stage_1_0_t352;
    FSM_dct_8x8_stage_1_0_t354 = FSM_dct_8x8_stage_1_0_t353[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t355 = FSM_dct_8x8_stage_1_0_t335;
    FSM_dct_8x8_stage_1_0_t355[FSM_dct_8x8_stage_1_0_t340 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t354;
    FSM_dct_8x8_stage_1_0_t356 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_1_0_t357 = FSM_dct_8x8_stage_1_0_t356[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t358 = FSM_dct_8x8_stage_1_0_t357 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_1_0_t359 = FSM_dct_8x8_stage_1_0_t358[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t360 = FSM_dct_8x8_stage_1_0_t359[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t361 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_1_0_t362 = FSM_dct_8x8_stage_1_0_t361[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t363 = FSM_dct_8x8_stage_1_0_t362 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_1_0_t364 = FSM_dct_8x8_stage_1_0_t363[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t365 = FSM_dct_8x8_stage_1_0_t364[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t366 = i_data_in[FSM_dct_8x8_stage_1_0_t365 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t367 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_1_0_t368 = FSM_dct_8x8_stage_1_0_t367[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t369 = FSM_dct_8x8_stage_1_0_t368 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_1_0_t370 = FSM_dct_8x8_stage_1_0_t369[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t371 = FSM_dct_8x8_stage_1_0_t370[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t372 = i_data_in[FSM_dct_8x8_stage_1_0_t371 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t373 = FSM_dct_8x8_stage_1_0_t366 + FSM_dct_8x8_stage_1_0_t372;
    FSM_dct_8x8_stage_1_0_t374 = FSM_dct_8x8_stage_1_0_t373[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t375 = FSM_dct_8x8_stage_1_0_t355;
    FSM_dct_8x8_stage_1_0_t375[FSM_dct_8x8_stage_1_0_t360 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t374;
    FSM_dct_8x8_stage_1_0_t376 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_1_0_t377 = FSM_dct_8x8_stage_1_0_t376[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t378 = FSM_dct_8x8_stage_1_0_t377 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_1_0_t379 = FSM_dct_8x8_stage_1_0_t378[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t380 = FSM_dct_8x8_stage_1_0_t379[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t381 = FSM_dct_8x8_stage_1_0_t375;
    FSM_dct_8x8_stage_1_0_t381[FSM_dct_8x8_stage_1_0_t380 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t366 - FSM_dct_8x8_stage_1_0_t372;
    FSM_dct_8x8_stage_1_0_t382 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_1_0_t383 = FSM_dct_8x8_stage_1_0_t382[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t384 = FSM_dct_8x8_stage_1_0_t383 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_1_0_t385 = FSM_dct_8x8_stage_1_0_t384[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t386 = FSM_dct_8x8_stage_1_0_t385[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t387 = FSM_dct_8x8_stage_1_0_t381;
    FSM_dct_8x8_stage_1_0_t387[FSM_dct_8x8_stage_1_0_t386 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t346 - FSM_dct_8x8_stage_1_0_t352;
    FSM_dct_8x8_stage_1_0_t388 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_1_0_t389 = FSM_dct_8x8_stage_1_0_t388[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t390 = FSM_dct_8x8_stage_1_0_t389 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_1_0_t391 = FSM_dct_8x8_stage_1_0_t390[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t392 = FSM_dct_8x8_stage_1_0_t391[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t393 = FSM_dct_8x8_stage_1_0_t387;
    FSM_dct_8x8_stage_1_0_t393[FSM_dct_8x8_stage_1_0_t392 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t326 - FSM_dct_8x8_stage_1_0_t332;
    FSM_dct_8x8_stage_1_0_t394 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_1_0_t395 = FSM_dct_8x8_stage_1_0_t394[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t396 = FSM_dct_8x8_stage_1_0_t395 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_1_0_t397 = FSM_dct_8x8_stage_1_0_t396[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t398 = FSM_dct_8x8_stage_1_0_t397[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t399 = FSM_dct_8x8_stage_1_0_t393;
    FSM_dct_8x8_stage_1_0_t399[FSM_dct_8x8_stage_1_0_t398 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t306 - FSM_dct_8x8_stage_1_0_t312;
    FSM_dct_8x8_stage_1_0_t400 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_1_0_t401 = FSM_dct_8x8_stage_1_0_t400[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t402 = FSM_dct_8x8_stage_1_0_t401[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t403 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_1_0_t404 = FSM_dct_8x8_stage_1_0_t403[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t405 = FSM_dct_8x8_stage_1_0_t404[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t406 = i_data_in[FSM_dct_8x8_stage_1_0_t405 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t407 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_1_0_t408 = FSM_dct_8x8_stage_1_0_t407[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t409 = FSM_dct_8x8_stage_1_0_t408 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_1_0_t410 = FSM_dct_8x8_stage_1_0_t409[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t411 = FSM_dct_8x8_stage_1_0_t410[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t412 = i_data_in[FSM_dct_8x8_stage_1_0_t411 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t413 = FSM_dct_8x8_stage_1_0_t406 + FSM_dct_8x8_stage_1_0_t412;
    FSM_dct_8x8_stage_1_0_t414 = FSM_dct_8x8_stage_1_0_t413[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t415 = FSM_dct_8x8_stage_1_0_t399;
    FSM_dct_8x8_stage_1_0_t415[FSM_dct_8x8_stage_1_0_t402 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t414;
    FSM_dct_8x8_stage_1_0_t416 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_1_0_t417 = FSM_dct_8x8_stage_1_0_t416[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t418 = FSM_dct_8x8_stage_1_0_t417 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_1_0_t419 = FSM_dct_8x8_stage_1_0_t418[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t420 = FSM_dct_8x8_stage_1_0_t419[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t421 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_1_0_t422 = FSM_dct_8x8_stage_1_0_t421[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t423 = FSM_dct_8x8_stage_1_0_t422 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_1_0_t424 = FSM_dct_8x8_stage_1_0_t423[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t425 = FSM_dct_8x8_stage_1_0_t424[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t426 = i_data_in[FSM_dct_8x8_stage_1_0_t425 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t427 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_1_0_t428 = FSM_dct_8x8_stage_1_0_t427[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t429 = FSM_dct_8x8_stage_1_0_t428 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_1_0_t430 = FSM_dct_8x8_stage_1_0_t429[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t431 = FSM_dct_8x8_stage_1_0_t430[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t432 = i_data_in[FSM_dct_8x8_stage_1_0_t431 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t433 = FSM_dct_8x8_stage_1_0_t426 + FSM_dct_8x8_stage_1_0_t432;
    FSM_dct_8x8_stage_1_0_t434 = FSM_dct_8x8_stage_1_0_t433[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t435 = FSM_dct_8x8_stage_1_0_t415;
    FSM_dct_8x8_stage_1_0_t435[FSM_dct_8x8_stage_1_0_t420 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t434;
    FSM_dct_8x8_stage_1_0_t436 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_1_0_t437 = FSM_dct_8x8_stage_1_0_t436[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t438 = FSM_dct_8x8_stage_1_0_t437 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_1_0_t439 = FSM_dct_8x8_stage_1_0_t438[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t440 = FSM_dct_8x8_stage_1_0_t439[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t441 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_1_0_t442 = FSM_dct_8x8_stage_1_0_t441[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t443 = FSM_dct_8x8_stage_1_0_t442 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_1_0_t444 = FSM_dct_8x8_stage_1_0_t443[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t445 = FSM_dct_8x8_stage_1_0_t444[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t446 = i_data_in[FSM_dct_8x8_stage_1_0_t445 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t447 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_1_0_t448 = FSM_dct_8x8_stage_1_0_t447[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t449 = FSM_dct_8x8_stage_1_0_t448 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_1_0_t450 = FSM_dct_8x8_stage_1_0_t449[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t451 = FSM_dct_8x8_stage_1_0_t450[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t452 = i_data_in[FSM_dct_8x8_stage_1_0_t451 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t453 = FSM_dct_8x8_stage_1_0_t446 + FSM_dct_8x8_stage_1_0_t452;
    FSM_dct_8x8_stage_1_0_t454 = FSM_dct_8x8_stage_1_0_t453[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t455 = FSM_dct_8x8_stage_1_0_t435;
    FSM_dct_8x8_stage_1_0_t455[FSM_dct_8x8_stage_1_0_t440 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t454;
    FSM_dct_8x8_stage_1_0_t456 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_1_0_t457 = FSM_dct_8x8_stage_1_0_t456[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t458 = FSM_dct_8x8_stage_1_0_t457 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_1_0_t459 = FSM_dct_8x8_stage_1_0_t458[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t460 = FSM_dct_8x8_stage_1_0_t459[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t461 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_1_0_t462 = FSM_dct_8x8_stage_1_0_t461[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t463 = FSM_dct_8x8_stage_1_0_t462 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_1_0_t464 = FSM_dct_8x8_stage_1_0_t463[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t465 = FSM_dct_8x8_stage_1_0_t464[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t466 = i_data_in[FSM_dct_8x8_stage_1_0_t465 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t467 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_1_0_t468 = FSM_dct_8x8_stage_1_0_t467[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t469 = FSM_dct_8x8_stage_1_0_t468 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_1_0_t470 = FSM_dct_8x8_stage_1_0_t469[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t471 = FSM_dct_8x8_stage_1_0_t470[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t472 = i_data_in[FSM_dct_8x8_stage_1_0_t471 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t473 = FSM_dct_8x8_stage_1_0_t466 + FSM_dct_8x8_stage_1_0_t472;
    FSM_dct_8x8_stage_1_0_t474 = FSM_dct_8x8_stage_1_0_t473[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t475 = FSM_dct_8x8_stage_1_0_t455;
    FSM_dct_8x8_stage_1_0_t475[FSM_dct_8x8_stage_1_0_t460 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t474;
    FSM_dct_8x8_stage_1_0_t476 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_1_0_t477 = FSM_dct_8x8_stage_1_0_t476[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t478 = FSM_dct_8x8_stage_1_0_t477 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_1_0_t479 = FSM_dct_8x8_stage_1_0_t478[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t480 = FSM_dct_8x8_stage_1_0_t479[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t481 = FSM_dct_8x8_stage_1_0_t475;
    FSM_dct_8x8_stage_1_0_t481[FSM_dct_8x8_stage_1_0_t480 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t466 - FSM_dct_8x8_stage_1_0_t472;
    FSM_dct_8x8_stage_1_0_t482 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_1_0_t483 = FSM_dct_8x8_stage_1_0_t482[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t484 = FSM_dct_8x8_stage_1_0_t483 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_1_0_t485 = FSM_dct_8x8_stage_1_0_t484[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t486 = FSM_dct_8x8_stage_1_0_t485[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t487 = FSM_dct_8x8_stage_1_0_t481;
    FSM_dct_8x8_stage_1_0_t487[FSM_dct_8x8_stage_1_0_t486 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t446 - FSM_dct_8x8_stage_1_0_t452;
    FSM_dct_8x8_stage_1_0_t488 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_1_0_t489 = FSM_dct_8x8_stage_1_0_t488[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t490 = FSM_dct_8x8_stage_1_0_t489 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_1_0_t491 = FSM_dct_8x8_stage_1_0_t490[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t492 = FSM_dct_8x8_stage_1_0_t491[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t493 = FSM_dct_8x8_stage_1_0_t487;
    FSM_dct_8x8_stage_1_0_t493[FSM_dct_8x8_stage_1_0_t492 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t426 - FSM_dct_8x8_stage_1_0_t432;
    FSM_dct_8x8_stage_1_0_t494 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_1_0_t495 = FSM_dct_8x8_stage_1_0_t494[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t496 = FSM_dct_8x8_stage_1_0_t495 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_1_0_t497 = FSM_dct_8x8_stage_1_0_t496[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t498 = FSM_dct_8x8_stage_1_0_t497[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t499 = FSM_dct_8x8_stage_1_0_t493;
    FSM_dct_8x8_stage_1_0_t499[FSM_dct_8x8_stage_1_0_t498 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t406 - FSM_dct_8x8_stage_1_0_t412;
    FSM_dct_8x8_stage_1_0_t500 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_1_0_t501 = FSM_dct_8x8_stage_1_0_t500[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t502 = FSM_dct_8x8_stage_1_0_t501[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t503 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_1_0_t504 = FSM_dct_8x8_stage_1_0_t503[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t505 = FSM_dct_8x8_stage_1_0_t504[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t506 = i_data_in[FSM_dct_8x8_stage_1_0_t505 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t507 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_1_0_t508 = FSM_dct_8x8_stage_1_0_t507[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t509 = FSM_dct_8x8_stage_1_0_t508 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_1_0_t510 = FSM_dct_8x8_stage_1_0_t509[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t511 = FSM_dct_8x8_stage_1_0_t510[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t512 = i_data_in[FSM_dct_8x8_stage_1_0_t511 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t513 = FSM_dct_8x8_stage_1_0_t506 + FSM_dct_8x8_stage_1_0_t512;
    FSM_dct_8x8_stage_1_0_t514 = FSM_dct_8x8_stage_1_0_t513[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t515 = FSM_dct_8x8_stage_1_0_t499;
    FSM_dct_8x8_stage_1_0_t515[FSM_dct_8x8_stage_1_0_t502 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t514;
    FSM_dct_8x8_stage_1_0_t516 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_1_0_t517 = FSM_dct_8x8_stage_1_0_t516[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t518 = FSM_dct_8x8_stage_1_0_t517 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_1_0_t519 = FSM_dct_8x8_stage_1_0_t518[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t520 = FSM_dct_8x8_stage_1_0_t519[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t521 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_1_0_t522 = FSM_dct_8x8_stage_1_0_t521[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t523 = FSM_dct_8x8_stage_1_0_t522 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_1_0_t524 = FSM_dct_8x8_stage_1_0_t523[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t525 = FSM_dct_8x8_stage_1_0_t524[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t526 = i_data_in[FSM_dct_8x8_stage_1_0_t525 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t527 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_1_0_t528 = FSM_dct_8x8_stage_1_0_t527[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t529 = FSM_dct_8x8_stage_1_0_t528 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_1_0_t530 = FSM_dct_8x8_stage_1_0_t529[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t531 = FSM_dct_8x8_stage_1_0_t530[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t532 = i_data_in[FSM_dct_8x8_stage_1_0_t531 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t533 = FSM_dct_8x8_stage_1_0_t526 + FSM_dct_8x8_stage_1_0_t532;
    FSM_dct_8x8_stage_1_0_t534 = FSM_dct_8x8_stage_1_0_t533[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t535 = FSM_dct_8x8_stage_1_0_t515;
    FSM_dct_8x8_stage_1_0_t535[FSM_dct_8x8_stage_1_0_t520 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t534;
    FSM_dct_8x8_stage_1_0_t536 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_1_0_t537 = FSM_dct_8x8_stage_1_0_t536[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t538 = FSM_dct_8x8_stage_1_0_t537 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_1_0_t539 = FSM_dct_8x8_stage_1_0_t538[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t540 = FSM_dct_8x8_stage_1_0_t539[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t541 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_1_0_t542 = FSM_dct_8x8_stage_1_0_t541[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t543 = FSM_dct_8x8_stage_1_0_t542 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_1_0_t544 = FSM_dct_8x8_stage_1_0_t543[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t545 = FSM_dct_8x8_stage_1_0_t544[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t546 = i_data_in[FSM_dct_8x8_stage_1_0_t545 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t547 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_1_0_t548 = FSM_dct_8x8_stage_1_0_t547[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t549 = FSM_dct_8x8_stage_1_0_t548 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_1_0_t550 = FSM_dct_8x8_stage_1_0_t549[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t551 = FSM_dct_8x8_stage_1_0_t550[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t552 = i_data_in[FSM_dct_8x8_stage_1_0_t551 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t553 = FSM_dct_8x8_stage_1_0_t546 + FSM_dct_8x8_stage_1_0_t552;
    FSM_dct_8x8_stage_1_0_t554 = FSM_dct_8x8_stage_1_0_t553[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t555 = FSM_dct_8x8_stage_1_0_t535;
    FSM_dct_8x8_stage_1_0_t555[FSM_dct_8x8_stage_1_0_t540 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t554;
    FSM_dct_8x8_stage_1_0_t556 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_1_0_t557 = FSM_dct_8x8_stage_1_0_t556[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t558 = FSM_dct_8x8_stage_1_0_t557 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_1_0_t559 = FSM_dct_8x8_stage_1_0_t558[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t560 = FSM_dct_8x8_stage_1_0_t559[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t561 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_1_0_t562 = FSM_dct_8x8_stage_1_0_t561[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t563 = FSM_dct_8x8_stage_1_0_t562 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_1_0_t564 = FSM_dct_8x8_stage_1_0_t563[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t565 = FSM_dct_8x8_stage_1_0_t564[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t566 = i_data_in[FSM_dct_8x8_stage_1_0_t565 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t567 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_1_0_t568 = FSM_dct_8x8_stage_1_0_t567[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t569 = FSM_dct_8x8_stage_1_0_t568 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_1_0_t570 = FSM_dct_8x8_stage_1_0_t569[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t571 = FSM_dct_8x8_stage_1_0_t570[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t572 = i_data_in[FSM_dct_8x8_stage_1_0_t571 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t573 = FSM_dct_8x8_stage_1_0_t566 + FSM_dct_8x8_stage_1_0_t572;
    FSM_dct_8x8_stage_1_0_t574 = FSM_dct_8x8_stage_1_0_t573[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t575 = FSM_dct_8x8_stage_1_0_t555;
    FSM_dct_8x8_stage_1_0_t575[FSM_dct_8x8_stage_1_0_t560 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t574;
    FSM_dct_8x8_stage_1_0_t576 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_1_0_t577 = FSM_dct_8x8_stage_1_0_t576[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t578 = FSM_dct_8x8_stage_1_0_t577 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_1_0_t579 = FSM_dct_8x8_stage_1_0_t578[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t580 = FSM_dct_8x8_stage_1_0_t579[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t581 = FSM_dct_8x8_stage_1_0_t575;
    FSM_dct_8x8_stage_1_0_t581[FSM_dct_8x8_stage_1_0_t580 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t566 - FSM_dct_8x8_stage_1_0_t572;
    FSM_dct_8x8_stage_1_0_t582 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_1_0_t583 = FSM_dct_8x8_stage_1_0_t582[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t584 = FSM_dct_8x8_stage_1_0_t583 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_1_0_t585 = FSM_dct_8x8_stage_1_0_t584[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t586 = FSM_dct_8x8_stage_1_0_t585[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t587 = FSM_dct_8x8_stage_1_0_t581;
    FSM_dct_8x8_stage_1_0_t587[FSM_dct_8x8_stage_1_0_t586 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t546 - FSM_dct_8x8_stage_1_0_t552;
    FSM_dct_8x8_stage_1_0_t588 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_1_0_t589 = FSM_dct_8x8_stage_1_0_t588[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t590 = FSM_dct_8x8_stage_1_0_t589 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_1_0_t591 = FSM_dct_8x8_stage_1_0_t590[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t592 = FSM_dct_8x8_stage_1_0_t591[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t593 = FSM_dct_8x8_stage_1_0_t587;
    FSM_dct_8x8_stage_1_0_t593[FSM_dct_8x8_stage_1_0_t592 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t526 - FSM_dct_8x8_stage_1_0_t532;
    FSM_dct_8x8_stage_1_0_t594 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_1_0_t595 = FSM_dct_8x8_stage_1_0_t594[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t596 = FSM_dct_8x8_stage_1_0_t595 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_1_0_t597 = FSM_dct_8x8_stage_1_0_t596[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t598 = FSM_dct_8x8_stage_1_0_t597[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t599 = FSM_dct_8x8_stage_1_0_t593;
    FSM_dct_8x8_stage_1_0_t599[FSM_dct_8x8_stage_1_0_t598 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t506 - FSM_dct_8x8_stage_1_0_t512;
    FSM_dct_8x8_stage_1_0_t600 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_1_0_t601 = FSM_dct_8x8_stage_1_0_t600[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t602 = FSM_dct_8x8_stage_1_0_t601[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t603 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_1_0_t604 = FSM_dct_8x8_stage_1_0_t603[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t605 = FSM_dct_8x8_stage_1_0_t604[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t606 = i_data_in[FSM_dct_8x8_stage_1_0_t605 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t607 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_1_0_t608 = FSM_dct_8x8_stage_1_0_t607[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t609 = FSM_dct_8x8_stage_1_0_t608 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_1_0_t610 = FSM_dct_8x8_stage_1_0_t609[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t611 = FSM_dct_8x8_stage_1_0_t610[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t612 = i_data_in[FSM_dct_8x8_stage_1_0_t611 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t613 = FSM_dct_8x8_stage_1_0_t606 + FSM_dct_8x8_stage_1_0_t612;
    FSM_dct_8x8_stage_1_0_t614 = FSM_dct_8x8_stage_1_0_t613[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t615 = FSM_dct_8x8_stage_1_0_t599;
    FSM_dct_8x8_stage_1_0_t615[FSM_dct_8x8_stage_1_0_t602 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t614;
    FSM_dct_8x8_stage_1_0_t616 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_1_0_t617 = FSM_dct_8x8_stage_1_0_t616[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t618 = FSM_dct_8x8_stage_1_0_t617 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_1_0_t619 = FSM_dct_8x8_stage_1_0_t618[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t620 = FSM_dct_8x8_stage_1_0_t619[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t621 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_1_0_t622 = FSM_dct_8x8_stage_1_0_t621[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t623 = FSM_dct_8x8_stage_1_0_t622 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_1_0_t624 = FSM_dct_8x8_stage_1_0_t623[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t625 = FSM_dct_8x8_stage_1_0_t624[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t626 = i_data_in[FSM_dct_8x8_stage_1_0_t625 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t627 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_1_0_t628 = FSM_dct_8x8_stage_1_0_t627[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t629 = FSM_dct_8x8_stage_1_0_t628 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_1_0_t630 = FSM_dct_8x8_stage_1_0_t629[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t631 = FSM_dct_8x8_stage_1_0_t630[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t632 = i_data_in[FSM_dct_8x8_stage_1_0_t631 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t633 = FSM_dct_8x8_stage_1_0_t626 + FSM_dct_8x8_stage_1_0_t632;
    FSM_dct_8x8_stage_1_0_t634 = FSM_dct_8x8_stage_1_0_t633[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t635 = FSM_dct_8x8_stage_1_0_t615;
    FSM_dct_8x8_stage_1_0_t635[FSM_dct_8x8_stage_1_0_t620 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t634;
    FSM_dct_8x8_stage_1_0_t636 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_1_0_t637 = FSM_dct_8x8_stage_1_0_t636[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t638 = FSM_dct_8x8_stage_1_0_t637 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_1_0_t639 = FSM_dct_8x8_stage_1_0_t638[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t640 = FSM_dct_8x8_stage_1_0_t639[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t641 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_1_0_t642 = FSM_dct_8x8_stage_1_0_t641[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t643 = FSM_dct_8x8_stage_1_0_t642 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_1_0_t644 = FSM_dct_8x8_stage_1_0_t643[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t645 = FSM_dct_8x8_stage_1_0_t644[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t646 = i_data_in[FSM_dct_8x8_stage_1_0_t645 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t647 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_1_0_t648 = FSM_dct_8x8_stage_1_0_t647[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t649 = FSM_dct_8x8_stage_1_0_t648 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_1_0_t650 = FSM_dct_8x8_stage_1_0_t649[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t651 = FSM_dct_8x8_stage_1_0_t650[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t652 = i_data_in[FSM_dct_8x8_stage_1_0_t651 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t653 = FSM_dct_8x8_stage_1_0_t646 + FSM_dct_8x8_stage_1_0_t652;
    FSM_dct_8x8_stage_1_0_t654 = FSM_dct_8x8_stage_1_0_t653[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t655 = FSM_dct_8x8_stage_1_0_t635;
    FSM_dct_8x8_stage_1_0_t655[FSM_dct_8x8_stage_1_0_t640 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t654;
    FSM_dct_8x8_stage_1_0_t656 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_1_0_t657 = FSM_dct_8x8_stage_1_0_t656[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t658 = FSM_dct_8x8_stage_1_0_t657 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_1_0_t659 = FSM_dct_8x8_stage_1_0_t658[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t660 = FSM_dct_8x8_stage_1_0_t659[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t661 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_1_0_t662 = FSM_dct_8x8_stage_1_0_t661[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t663 = FSM_dct_8x8_stage_1_0_t662 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_1_0_t664 = FSM_dct_8x8_stage_1_0_t663[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t665 = FSM_dct_8x8_stage_1_0_t664[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t666 = i_data_in[FSM_dct_8x8_stage_1_0_t665 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t667 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_1_0_t668 = FSM_dct_8x8_stage_1_0_t667[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t669 = FSM_dct_8x8_stage_1_0_t668 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_1_0_t670 = FSM_dct_8x8_stage_1_0_t669[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t671 = FSM_dct_8x8_stage_1_0_t670[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t672 = i_data_in[FSM_dct_8x8_stage_1_0_t671 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t673 = FSM_dct_8x8_stage_1_0_t666 + FSM_dct_8x8_stage_1_0_t672;
    FSM_dct_8x8_stage_1_0_t674 = FSM_dct_8x8_stage_1_0_t673[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t675 = FSM_dct_8x8_stage_1_0_t655;
    FSM_dct_8x8_stage_1_0_t675[FSM_dct_8x8_stage_1_0_t660 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t674;
    FSM_dct_8x8_stage_1_0_t676 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_1_0_t677 = FSM_dct_8x8_stage_1_0_t676[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t678 = FSM_dct_8x8_stage_1_0_t677 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_1_0_t679 = FSM_dct_8x8_stage_1_0_t678[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t680 = FSM_dct_8x8_stage_1_0_t679[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t681 = FSM_dct_8x8_stage_1_0_t675;
    FSM_dct_8x8_stage_1_0_t681[FSM_dct_8x8_stage_1_0_t680 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t666 - FSM_dct_8x8_stage_1_0_t672;
    FSM_dct_8x8_stage_1_0_t682 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_1_0_t683 = FSM_dct_8x8_stage_1_0_t682[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t684 = FSM_dct_8x8_stage_1_0_t683 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_1_0_t685 = FSM_dct_8x8_stage_1_0_t684[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t686 = FSM_dct_8x8_stage_1_0_t685[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t687 = FSM_dct_8x8_stage_1_0_t681;
    FSM_dct_8x8_stage_1_0_t687[FSM_dct_8x8_stage_1_0_t686 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t646 - FSM_dct_8x8_stage_1_0_t652;
    FSM_dct_8x8_stage_1_0_t688 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_1_0_t689 = FSM_dct_8x8_stage_1_0_t688[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t690 = FSM_dct_8x8_stage_1_0_t689 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_1_0_t691 = FSM_dct_8x8_stage_1_0_t690[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t692 = FSM_dct_8x8_stage_1_0_t691[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t693 = FSM_dct_8x8_stage_1_0_t687;
    FSM_dct_8x8_stage_1_0_t693[FSM_dct_8x8_stage_1_0_t692 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t626 - FSM_dct_8x8_stage_1_0_t632;
    FSM_dct_8x8_stage_1_0_t694 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_1_0_t695 = FSM_dct_8x8_stage_1_0_t694[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t696 = FSM_dct_8x8_stage_1_0_t695 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_1_0_t697 = FSM_dct_8x8_stage_1_0_t696[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t698 = FSM_dct_8x8_stage_1_0_t697[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t699 = FSM_dct_8x8_stage_1_0_t693;
    FSM_dct_8x8_stage_1_0_t699[FSM_dct_8x8_stage_1_0_t698 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t606 - FSM_dct_8x8_stage_1_0_t612;
    FSM_dct_8x8_stage_1_0_t700 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_1_0_t701 = FSM_dct_8x8_stage_1_0_t700[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t702 = FSM_dct_8x8_stage_1_0_t701[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t703 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_1_0_t704 = FSM_dct_8x8_stage_1_0_t703[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t705 = FSM_dct_8x8_stage_1_0_t704[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t706 = i_data_in[FSM_dct_8x8_stage_1_0_t705 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t707 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_1_0_t708 = FSM_dct_8x8_stage_1_0_t707[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t709 = FSM_dct_8x8_stage_1_0_t708 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_1_0_t710 = FSM_dct_8x8_stage_1_0_t709[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t711 = FSM_dct_8x8_stage_1_0_t710[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t712 = i_data_in[FSM_dct_8x8_stage_1_0_t711 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t713 = FSM_dct_8x8_stage_1_0_t706 + FSM_dct_8x8_stage_1_0_t712;
    FSM_dct_8x8_stage_1_0_t714 = FSM_dct_8x8_stage_1_0_t713[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t715 = FSM_dct_8x8_stage_1_0_t699;
    FSM_dct_8x8_stage_1_0_t715[FSM_dct_8x8_stage_1_0_t702 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t714;
    FSM_dct_8x8_stage_1_0_t716 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_1_0_t717 = FSM_dct_8x8_stage_1_0_t716[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t718 = FSM_dct_8x8_stage_1_0_t717 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_1_0_t719 = FSM_dct_8x8_stage_1_0_t718[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t720 = FSM_dct_8x8_stage_1_0_t719[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t721 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_1_0_t722 = FSM_dct_8x8_stage_1_0_t721[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t723 = FSM_dct_8x8_stage_1_0_t722 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_1_0_t724 = FSM_dct_8x8_stage_1_0_t723[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t725 = FSM_dct_8x8_stage_1_0_t724[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t726 = i_data_in[FSM_dct_8x8_stage_1_0_t725 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t727 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_1_0_t728 = FSM_dct_8x8_stage_1_0_t727[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t729 = FSM_dct_8x8_stage_1_0_t728 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_1_0_t730 = FSM_dct_8x8_stage_1_0_t729[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t731 = FSM_dct_8x8_stage_1_0_t730[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t732 = i_data_in[FSM_dct_8x8_stage_1_0_t731 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t733 = FSM_dct_8x8_stage_1_0_t726 + FSM_dct_8x8_stage_1_0_t732;
    FSM_dct_8x8_stage_1_0_t734 = FSM_dct_8x8_stage_1_0_t733[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t735 = FSM_dct_8x8_stage_1_0_t715;
    FSM_dct_8x8_stage_1_0_t735[FSM_dct_8x8_stage_1_0_t720 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t734;
    FSM_dct_8x8_stage_1_0_t736 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_1_0_t737 = FSM_dct_8x8_stage_1_0_t736[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t738 = FSM_dct_8x8_stage_1_0_t737 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_1_0_t739 = FSM_dct_8x8_stage_1_0_t738[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t740 = FSM_dct_8x8_stage_1_0_t739[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t741 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_1_0_t742 = FSM_dct_8x8_stage_1_0_t741[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t743 = FSM_dct_8x8_stage_1_0_t742 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_1_0_t744 = FSM_dct_8x8_stage_1_0_t743[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t745 = FSM_dct_8x8_stage_1_0_t744[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t746 = i_data_in[FSM_dct_8x8_stage_1_0_t745 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t747 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_1_0_t748 = FSM_dct_8x8_stage_1_0_t747[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t749 = FSM_dct_8x8_stage_1_0_t748 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_1_0_t750 = FSM_dct_8x8_stage_1_0_t749[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t751 = FSM_dct_8x8_stage_1_0_t750[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t752 = i_data_in[FSM_dct_8x8_stage_1_0_t751 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t753 = FSM_dct_8x8_stage_1_0_t746 + FSM_dct_8x8_stage_1_0_t752;
    FSM_dct_8x8_stage_1_0_t754 = FSM_dct_8x8_stage_1_0_t753[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t755 = FSM_dct_8x8_stage_1_0_t735;
    FSM_dct_8x8_stage_1_0_t755[FSM_dct_8x8_stage_1_0_t740 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t754;
    FSM_dct_8x8_stage_1_0_t756 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_1_0_t757 = FSM_dct_8x8_stage_1_0_t756[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t758 = FSM_dct_8x8_stage_1_0_t757 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_1_0_t759 = FSM_dct_8x8_stage_1_0_t758[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t760 = FSM_dct_8x8_stage_1_0_t759[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t761 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_1_0_t762 = FSM_dct_8x8_stage_1_0_t761[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t763 = FSM_dct_8x8_stage_1_0_t762 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_1_0_t764 = FSM_dct_8x8_stage_1_0_t763[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t765 = FSM_dct_8x8_stage_1_0_t764[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t766 = i_data_in[FSM_dct_8x8_stage_1_0_t765 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t767 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_1_0_t768 = FSM_dct_8x8_stage_1_0_t767[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t769 = FSM_dct_8x8_stage_1_0_t768 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_1_0_t770 = FSM_dct_8x8_stage_1_0_t769[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t771 = FSM_dct_8x8_stage_1_0_t770[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t772 = i_data_in[FSM_dct_8x8_stage_1_0_t771 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t773 = FSM_dct_8x8_stage_1_0_t766 + FSM_dct_8x8_stage_1_0_t772;
    FSM_dct_8x8_stage_1_0_t774 = FSM_dct_8x8_stage_1_0_t773[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t775 = FSM_dct_8x8_stage_1_0_t755;
    FSM_dct_8x8_stage_1_0_t775[FSM_dct_8x8_stage_1_0_t760 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t774;
    FSM_dct_8x8_stage_1_0_t776 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_1_0_t777 = FSM_dct_8x8_stage_1_0_t776[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t778 = FSM_dct_8x8_stage_1_0_t777 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_1_0_t779 = FSM_dct_8x8_stage_1_0_t778[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t780 = FSM_dct_8x8_stage_1_0_t779[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t781 = FSM_dct_8x8_stage_1_0_t775;
    FSM_dct_8x8_stage_1_0_t781[FSM_dct_8x8_stage_1_0_t780 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t766 - FSM_dct_8x8_stage_1_0_t772;
    FSM_dct_8x8_stage_1_0_t782 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_1_0_t783 = FSM_dct_8x8_stage_1_0_t782[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t784 = FSM_dct_8x8_stage_1_0_t783 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_1_0_t785 = FSM_dct_8x8_stage_1_0_t784[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t786 = FSM_dct_8x8_stage_1_0_t785[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t787 = FSM_dct_8x8_stage_1_0_t781;
    FSM_dct_8x8_stage_1_0_t787[FSM_dct_8x8_stage_1_0_t786 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t746 - FSM_dct_8x8_stage_1_0_t752;
    FSM_dct_8x8_stage_1_0_t788 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_1_0_t789 = FSM_dct_8x8_stage_1_0_t788[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t790 = FSM_dct_8x8_stage_1_0_t789 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_1_0_t791 = FSM_dct_8x8_stage_1_0_t790[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t792 = FSM_dct_8x8_stage_1_0_t791[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t793 = FSM_dct_8x8_stage_1_0_t787;
    FSM_dct_8x8_stage_1_0_t793[FSM_dct_8x8_stage_1_0_t792 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t726 - FSM_dct_8x8_stage_1_0_t732;
    FSM_dct_8x8_stage_1_0_t794 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_1_0_t795 = FSM_dct_8x8_stage_1_0_t794[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t796 = FSM_dct_8x8_stage_1_0_t795 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_1_0_t797 = FSM_dct_8x8_stage_1_0_t796[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t798 = FSM_dct_8x8_stage_1_0_t797[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t799 = FSM_dct_8x8_stage_1_0_t793;
    FSM_dct_8x8_stage_1_0_t799[FSM_dct_8x8_stage_1_0_t798 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t706 - FSM_dct_8x8_stage_1_0_t712;
end

always @* begin
    FSM_dct_8x8_stage_1_0_t0 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_1_0_t1 = FSM_dct_8x8_stage_1_0_t0[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t2 = FSM_dct_8x8_stage_1_0_t1[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t3 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_1_0_t4 = FSM_dct_8x8_stage_1_0_t3[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t5 = FSM_dct_8x8_stage_1_0_t4[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t6 = i_data_in[FSM_dct_8x8_stage_1_0_t5 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t7 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_1_0_t8 = FSM_dct_8x8_stage_1_0_t7[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t9 = FSM_dct_8x8_stage_1_0_t8 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_1_0_t10 = FSM_dct_8x8_stage_1_0_t9[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t11 = FSM_dct_8x8_stage_1_0_t10[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t12 = i_data_in[FSM_dct_8x8_stage_1_0_t11 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t13 = FSM_dct_8x8_stage_1_0_t6 + FSM_dct_8x8_stage_1_0_t12;
    FSM_dct_8x8_stage_1_0_t14 = FSM_dct_8x8_stage_1_0_t13[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t15 = 2048'b0;
    FSM_dct_8x8_stage_1_0_t15[FSM_dct_8x8_stage_1_0_t2 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t14;
    FSM_dct_8x8_stage_1_0_t16 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_1_0_t17 = FSM_dct_8x8_stage_1_0_t16[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t18 = FSM_dct_8x8_stage_1_0_t17 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_1_0_t19 = FSM_dct_8x8_stage_1_0_t18[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t20 = FSM_dct_8x8_stage_1_0_t19[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t21 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_1_0_t22 = FSM_dct_8x8_stage_1_0_t21[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t23 = FSM_dct_8x8_stage_1_0_t22 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_1_0_t24 = FSM_dct_8x8_stage_1_0_t23[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t25 = FSM_dct_8x8_stage_1_0_t24[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t26 = i_data_in[FSM_dct_8x8_stage_1_0_t25 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t27 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_1_0_t28 = FSM_dct_8x8_stage_1_0_t27[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t29 = FSM_dct_8x8_stage_1_0_t28 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_1_0_t30 = FSM_dct_8x8_stage_1_0_t29[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t31 = FSM_dct_8x8_stage_1_0_t30[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t32 = i_data_in[FSM_dct_8x8_stage_1_0_t31 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t33 = FSM_dct_8x8_stage_1_0_t26 + FSM_dct_8x8_stage_1_0_t32;
    FSM_dct_8x8_stage_1_0_t34 = FSM_dct_8x8_stage_1_0_t33[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t35 = FSM_dct_8x8_stage_1_0_t15;
    FSM_dct_8x8_stage_1_0_t35[FSM_dct_8x8_stage_1_0_t20 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t34;
    FSM_dct_8x8_stage_1_0_t36 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_1_0_t37 = FSM_dct_8x8_stage_1_0_t36[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t38 = FSM_dct_8x8_stage_1_0_t37 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_1_0_t39 = FSM_dct_8x8_stage_1_0_t38[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t40 = FSM_dct_8x8_stage_1_0_t39[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t41 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_1_0_t42 = FSM_dct_8x8_stage_1_0_t41[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t43 = FSM_dct_8x8_stage_1_0_t42 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_1_0_t44 = FSM_dct_8x8_stage_1_0_t43[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t45 = FSM_dct_8x8_stage_1_0_t44[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t46 = i_data_in[FSM_dct_8x8_stage_1_0_t45 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t47 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_1_0_t48 = FSM_dct_8x8_stage_1_0_t47[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t49 = FSM_dct_8x8_stage_1_0_t48 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_1_0_t50 = FSM_dct_8x8_stage_1_0_t49[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t51 = FSM_dct_8x8_stage_1_0_t50[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t52 = i_data_in[FSM_dct_8x8_stage_1_0_t51 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t53 = FSM_dct_8x8_stage_1_0_t46 + FSM_dct_8x8_stage_1_0_t52;
    FSM_dct_8x8_stage_1_0_t54 = FSM_dct_8x8_stage_1_0_t53[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t55 = FSM_dct_8x8_stage_1_0_t35;
    FSM_dct_8x8_stage_1_0_t55[FSM_dct_8x8_stage_1_0_t40 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t54;
    FSM_dct_8x8_stage_1_0_t56 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_1_0_t57 = FSM_dct_8x8_stage_1_0_t56[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t58 = FSM_dct_8x8_stage_1_0_t57 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_1_0_t59 = FSM_dct_8x8_stage_1_0_t58[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t60 = FSM_dct_8x8_stage_1_0_t59[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t61 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_1_0_t62 = FSM_dct_8x8_stage_1_0_t61[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t63 = FSM_dct_8x8_stage_1_0_t62 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_1_0_t64 = FSM_dct_8x8_stage_1_0_t63[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t65 = FSM_dct_8x8_stage_1_0_t64[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t66 = i_data_in[FSM_dct_8x8_stage_1_0_t65 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t67 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_1_0_t68 = FSM_dct_8x8_stage_1_0_t67[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t69 = FSM_dct_8x8_stage_1_0_t68 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_1_0_t70 = FSM_dct_8x8_stage_1_0_t69[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t71 = FSM_dct_8x8_stage_1_0_t70[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t72 = i_data_in[FSM_dct_8x8_stage_1_0_t71 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t73 = FSM_dct_8x8_stage_1_0_t66 + FSM_dct_8x8_stage_1_0_t72;
    FSM_dct_8x8_stage_1_0_t74 = FSM_dct_8x8_stage_1_0_t73[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t75 = FSM_dct_8x8_stage_1_0_t55;
    FSM_dct_8x8_stage_1_0_t75[FSM_dct_8x8_stage_1_0_t60 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t74;
    FSM_dct_8x8_stage_1_0_t76 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_1_0_t77 = FSM_dct_8x8_stage_1_0_t76[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t78 = FSM_dct_8x8_stage_1_0_t77 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_1_0_t79 = FSM_dct_8x8_stage_1_0_t78[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t80 = FSM_dct_8x8_stage_1_0_t79[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t81 = FSM_dct_8x8_stage_1_0_t75;
    FSM_dct_8x8_stage_1_0_t81[FSM_dct_8x8_stage_1_0_t80 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t66 - FSM_dct_8x8_stage_1_0_t72;
    FSM_dct_8x8_stage_1_0_t82 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_1_0_t83 = FSM_dct_8x8_stage_1_0_t82[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t84 = FSM_dct_8x8_stage_1_0_t83 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_1_0_t85 = FSM_dct_8x8_stage_1_0_t84[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t86 = FSM_dct_8x8_stage_1_0_t85[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t87 = FSM_dct_8x8_stage_1_0_t81;
    FSM_dct_8x8_stage_1_0_t87[FSM_dct_8x8_stage_1_0_t86 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t46 - FSM_dct_8x8_stage_1_0_t52;
    FSM_dct_8x8_stage_1_0_t88 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_1_0_t89 = FSM_dct_8x8_stage_1_0_t88[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t90 = FSM_dct_8x8_stage_1_0_t89 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_1_0_t91 = FSM_dct_8x8_stage_1_0_t90[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t92 = FSM_dct_8x8_stage_1_0_t91[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t93 = FSM_dct_8x8_stage_1_0_t87;
    FSM_dct_8x8_stage_1_0_t93[FSM_dct_8x8_stage_1_0_t92 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t26 - FSM_dct_8x8_stage_1_0_t32;
    FSM_dct_8x8_stage_1_0_t94 = 32'b00000000000000000000000000001000 * 32'b0;
    FSM_dct_8x8_stage_1_0_t95 = FSM_dct_8x8_stage_1_0_t94[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t96 = FSM_dct_8x8_stage_1_0_t95 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_1_0_t97 = FSM_dct_8x8_stage_1_0_t96[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t98 = FSM_dct_8x8_stage_1_0_t97[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t99 = FSM_dct_8x8_stage_1_0_t93;
    FSM_dct_8x8_stage_1_0_t99[FSM_dct_8x8_stage_1_0_t98 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t6 - FSM_dct_8x8_stage_1_0_t12;
    FSM_dct_8x8_stage_1_0_t100 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_1_0_t101 = FSM_dct_8x8_stage_1_0_t100[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t102 = FSM_dct_8x8_stage_1_0_t101[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t103 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_1_0_t104 = FSM_dct_8x8_stage_1_0_t103[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t105 = FSM_dct_8x8_stage_1_0_t104[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t106 = i_data_in[FSM_dct_8x8_stage_1_0_t105 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t107 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_1_0_t108 = FSM_dct_8x8_stage_1_0_t107[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t109 = FSM_dct_8x8_stage_1_0_t108 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_1_0_t110 = FSM_dct_8x8_stage_1_0_t109[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t111 = FSM_dct_8x8_stage_1_0_t110[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t112 = i_data_in[FSM_dct_8x8_stage_1_0_t111 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t113 = FSM_dct_8x8_stage_1_0_t106 + FSM_dct_8x8_stage_1_0_t112;
    FSM_dct_8x8_stage_1_0_t114 = FSM_dct_8x8_stage_1_0_t113[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t115 = FSM_dct_8x8_stage_1_0_t99;
    FSM_dct_8x8_stage_1_0_t115[FSM_dct_8x8_stage_1_0_t102 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t114;
    FSM_dct_8x8_stage_1_0_t116 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_1_0_t117 = FSM_dct_8x8_stage_1_0_t116[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t118 = FSM_dct_8x8_stage_1_0_t117 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_1_0_t119 = FSM_dct_8x8_stage_1_0_t118[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t120 = FSM_dct_8x8_stage_1_0_t119[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t121 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_1_0_t122 = FSM_dct_8x8_stage_1_0_t121[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t123 = FSM_dct_8x8_stage_1_0_t122 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_1_0_t124 = FSM_dct_8x8_stage_1_0_t123[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t125 = FSM_dct_8x8_stage_1_0_t124[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t126 = i_data_in[FSM_dct_8x8_stage_1_0_t125 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t127 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_1_0_t128 = FSM_dct_8x8_stage_1_0_t127[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t129 = FSM_dct_8x8_stage_1_0_t128 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_1_0_t130 = FSM_dct_8x8_stage_1_0_t129[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t131 = FSM_dct_8x8_stage_1_0_t130[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t132 = i_data_in[FSM_dct_8x8_stage_1_0_t131 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t133 = FSM_dct_8x8_stage_1_0_t126 + FSM_dct_8x8_stage_1_0_t132;
    FSM_dct_8x8_stage_1_0_t134 = FSM_dct_8x8_stage_1_0_t133[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t135 = FSM_dct_8x8_stage_1_0_t115;
    FSM_dct_8x8_stage_1_0_t135[FSM_dct_8x8_stage_1_0_t120 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t134;
    FSM_dct_8x8_stage_1_0_t136 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_1_0_t137 = FSM_dct_8x8_stage_1_0_t136[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t138 = FSM_dct_8x8_stage_1_0_t137 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_1_0_t139 = FSM_dct_8x8_stage_1_0_t138[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t140 = FSM_dct_8x8_stage_1_0_t139[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t141 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_1_0_t142 = FSM_dct_8x8_stage_1_0_t141[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t143 = FSM_dct_8x8_stage_1_0_t142 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_1_0_t144 = FSM_dct_8x8_stage_1_0_t143[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t145 = FSM_dct_8x8_stage_1_0_t144[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t146 = i_data_in[FSM_dct_8x8_stage_1_0_t145 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t147 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_1_0_t148 = FSM_dct_8x8_stage_1_0_t147[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t149 = FSM_dct_8x8_stage_1_0_t148 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_1_0_t150 = FSM_dct_8x8_stage_1_0_t149[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t151 = FSM_dct_8x8_stage_1_0_t150[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t152 = i_data_in[FSM_dct_8x8_stage_1_0_t151 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t153 = FSM_dct_8x8_stage_1_0_t146 + FSM_dct_8x8_stage_1_0_t152;
    FSM_dct_8x8_stage_1_0_t154 = FSM_dct_8x8_stage_1_0_t153[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t155 = FSM_dct_8x8_stage_1_0_t135;
    FSM_dct_8x8_stage_1_0_t155[FSM_dct_8x8_stage_1_0_t140 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t154;
    FSM_dct_8x8_stage_1_0_t156 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_1_0_t157 = FSM_dct_8x8_stage_1_0_t156[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t158 = FSM_dct_8x8_stage_1_0_t157 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_1_0_t159 = FSM_dct_8x8_stage_1_0_t158[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t160 = FSM_dct_8x8_stage_1_0_t159[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t161 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_1_0_t162 = FSM_dct_8x8_stage_1_0_t161[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t163 = FSM_dct_8x8_stage_1_0_t162 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_1_0_t164 = FSM_dct_8x8_stage_1_0_t163[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t165 = FSM_dct_8x8_stage_1_0_t164[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t166 = i_data_in[FSM_dct_8x8_stage_1_0_t165 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t167 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_1_0_t168 = FSM_dct_8x8_stage_1_0_t167[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t169 = FSM_dct_8x8_stage_1_0_t168 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_1_0_t170 = FSM_dct_8x8_stage_1_0_t169[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t171 = FSM_dct_8x8_stage_1_0_t170[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t172 = i_data_in[FSM_dct_8x8_stage_1_0_t171 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t173 = FSM_dct_8x8_stage_1_0_t166 + FSM_dct_8x8_stage_1_0_t172;
    FSM_dct_8x8_stage_1_0_t174 = FSM_dct_8x8_stage_1_0_t173[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t175 = FSM_dct_8x8_stage_1_0_t155;
    FSM_dct_8x8_stage_1_0_t175[FSM_dct_8x8_stage_1_0_t160 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t174;
    FSM_dct_8x8_stage_1_0_t176 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_1_0_t177 = FSM_dct_8x8_stage_1_0_t176[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t178 = FSM_dct_8x8_stage_1_0_t177 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_1_0_t179 = FSM_dct_8x8_stage_1_0_t178[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t180 = FSM_dct_8x8_stage_1_0_t179[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t181 = FSM_dct_8x8_stage_1_0_t175;
    FSM_dct_8x8_stage_1_0_t181[FSM_dct_8x8_stage_1_0_t180 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t166 - FSM_dct_8x8_stage_1_0_t172;
    FSM_dct_8x8_stage_1_0_t182 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_1_0_t183 = FSM_dct_8x8_stage_1_0_t182[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t184 = FSM_dct_8x8_stage_1_0_t183 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_1_0_t185 = FSM_dct_8x8_stage_1_0_t184[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t186 = FSM_dct_8x8_stage_1_0_t185[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t187 = FSM_dct_8x8_stage_1_0_t181;
    FSM_dct_8x8_stage_1_0_t187[FSM_dct_8x8_stage_1_0_t186 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t146 - FSM_dct_8x8_stage_1_0_t152;
    FSM_dct_8x8_stage_1_0_t188 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_1_0_t189 = FSM_dct_8x8_stage_1_0_t188[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t190 = FSM_dct_8x8_stage_1_0_t189 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_1_0_t191 = FSM_dct_8x8_stage_1_0_t190[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t192 = FSM_dct_8x8_stage_1_0_t191[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t193 = FSM_dct_8x8_stage_1_0_t187;
    FSM_dct_8x8_stage_1_0_t193[FSM_dct_8x8_stage_1_0_t192 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t126 - FSM_dct_8x8_stage_1_0_t132;
    FSM_dct_8x8_stage_1_0_t194 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_1_0_t195 = FSM_dct_8x8_stage_1_0_t194[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t196 = FSM_dct_8x8_stage_1_0_t195 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_1_0_t197 = FSM_dct_8x8_stage_1_0_t196[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t198 = FSM_dct_8x8_stage_1_0_t197[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t199 = FSM_dct_8x8_stage_1_0_t193;
    FSM_dct_8x8_stage_1_0_t199[FSM_dct_8x8_stage_1_0_t198 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t106 - FSM_dct_8x8_stage_1_0_t112;
    FSM_dct_8x8_stage_1_0_t200 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_1_0_t201 = FSM_dct_8x8_stage_1_0_t200[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t202 = FSM_dct_8x8_stage_1_0_t201[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t203 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_1_0_t204 = FSM_dct_8x8_stage_1_0_t203[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t205 = FSM_dct_8x8_stage_1_0_t204[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t206 = i_data_in[FSM_dct_8x8_stage_1_0_t205 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t207 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_1_0_t208 = FSM_dct_8x8_stage_1_0_t207[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t209 = FSM_dct_8x8_stage_1_0_t208 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_1_0_t210 = FSM_dct_8x8_stage_1_0_t209[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t211 = FSM_dct_8x8_stage_1_0_t210[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t212 = i_data_in[FSM_dct_8x8_stage_1_0_t211 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t213 = FSM_dct_8x8_stage_1_0_t206 + FSM_dct_8x8_stage_1_0_t212;
    FSM_dct_8x8_stage_1_0_t214 = FSM_dct_8x8_stage_1_0_t213[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t215 = FSM_dct_8x8_stage_1_0_t199;
    FSM_dct_8x8_stage_1_0_t215[FSM_dct_8x8_stage_1_0_t202 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t214;
    FSM_dct_8x8_stage_1_0_t216 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_1_0_t217 = FSM_dct_8x8_stage_1_0_t216[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t218 = FSM_dct_8x8_stage_1_0_t217 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_1_0_t219 = FSM_dct_8x8_stage_1_0_t218[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t220 = FSM_dct_8x8_stage_1_0_t219[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t221 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_1_0_t222 = FSM_dct_8x8_stage_1_0_t221[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t223 = FSM_dct_8x8_stage_1_0_t222 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_1_0_t224 = FSM_dct_8x8_stage_1_0_t223[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t225 = FSM_dct_8x8_stage_1_0_t224[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t226 = i_data_in[FSM_dct_8x8_stage_1_0_t225 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t227 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_1_0_t228 = FSM_dct_8x8_stage_1_0_t227[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t229 = FSM_dct_8x8_stage_1_0_t228 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_1_0_t230 = FSM_dct_8x8_stage_1_0_t229[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t231 = FSM_dct_8x8_stage_1_0_t230[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t232 = i_data_in[FSM_dct_8x8_stage_1_0_t231 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t233 = FSM_dct_8x8_stage_1_0_t226 + FSM_dct_8x8_stage_1_0_t232;
    FSM_dct_8x8_stage_1_0_t234 = FSM_dct_8x8_stage_1_0_t233[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t235 = FSM_dct_8x8_stage_1_0_t215;
    FSM_dct_8x8_stage_1_0_t235[FSM_dct_8x8_stage_1_0_t220 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t234;
    FSM_dct_8x8_stage_1_0_t236 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_1_0_t237 = FSM_dct_8x8_stage_1_0_t236[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t238 = FSM_dct_8x8_stage_1_0_t237 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_1_0_t239 = FSM_dct_8x8_stage_1_0_t238[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t240 = FSM_dct_8x8_stage_1_0_t239[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t241 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_1_0_t242 = FSM_dct_8x8_stage_1_0_t241[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t243 = FSM_dct_8x8_stage_1_0_t242 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_1_0_t244 = FSM_dct_8x8_stage_1_0_t243[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t245 = FSM_dct_8x8_stage_1_0_t244[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t246 = i_data_in[FSM_dct_8x8_stage_1_0_t245 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t247 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_1_0_t248 = FSM_dct_8x8_stage_1_0_t247[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t249 = FSM_dct_8x8_stage_1_0_t248 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_1_0_t250 = FSM_dct_8x8_stage_1_0_t249[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t251 = FSM_dct_8x8_stage_1_0_t250[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t252 = i_data_in[FSM_dct_8x8_stage_1_0_t251 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t253 = FSM_dct_8x8_stage_1_0_t246 + FSM_dct_8x8_stage_1_0_t252;
    FSM_dct_8x8_stage_1_0_t254 = FSM_dct_8x8_stage_1_0_t253[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t255 = FSM_dct_8x8_stage_1_0_t235;
    FSM_dct_8x8_stage_1_0_t255[FSM_dct_8x8_stage_1_0_t240 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t254;
    FSM_dct_8x8_stage_1_0_t256 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_1_0_t257 = FSM_dct_8x8_stage_1_0_t256[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t258 = FSM_dct_8x8_stage_1_0_t257 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_1_0_t259 = FSM_dct_8x8_stage_1_0_t258[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t260 = FSM_dct_8x8_stage_1_0_t259[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t261 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_1_0_t262 = FSM_dct_8x8_stage_1_0_t261[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t263 = FSM_dct_8x8_stage_1_0_t262 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_1_0_t264 = FSM_dct_8x8_stage_1_0_t263[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t265 = FSM_dct_8x8_stage_1_0_t264[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t266 = i_data_in[FSM_dct_8x8_stage_1_0_t265 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t267 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_1_0_t268 = FSM_dct_8x8_stage_1_0_t267[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t269 = FSM_dct_8x8_stage_1_0_t268 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_1_0_t270 = FSM_dct_8x8_stage_1_0_t269[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t271 = FSM_dct_8x8_stage_1_0_t270[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t272 = i_data_in[FSM_dct_8x8_stage_1_0_t271 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t273 = FSM_dct_8x8_stage_1_0_t266 + FSM_dct_8x8_stage_1_0_t272;
    FSM_dct_8x8_stage_1_0_t274 = FSM_dct_8x8_stage_1_0_t273[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t275 = FSM_dct_8x8_stage_1_0_t255;
    FSM_dct_8x8_stage_1_0_t275[FSM_dct_8x8_stage_1_0_t260 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t274;
    FSM_dct_8x8_stage_1_0_t276 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_1_0_t277 = FSM_dct_8x8_stage_1_0_t276[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t278 = FSM_dct_8x8_stage_1_0_t277 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_1_0_t279 = FSM_dct_8x8_stage_1_0_t278[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t280 = FSM_dct_8x8_stage_1_0_t279[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t281 = FSM_dct_8x8_stage_1_0_t275;
    FSM_dct_8x8_stage_1_0_t281[FSM_dct_8x8_stage_1_0_t280 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t266 - FSM_dct_8x8_stage_1_0_t272;
    FSM_dct_8x8_stage_1_0_t282 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_1_0_t283 = FSM_dct_8x8_stage_1_0_t282[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t284 = FSM_dct_8x8_stage_1_0_t283 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_1_0_t285 = FSM_dct_8x8_stage_1_0_t284[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t286 = FSM_dct_8x8_stage_1_0_t285[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t287 = FSM_dct_8x8_stage_1_0_t281;
    FSM_dct_8x8_stage_1_0_t287[FSM_dct_8x8_stage_1_0_t286 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t246 - FSM_dct_8x8_stage_1_0_t252;
    FSM_dct_8x8_stage_1_0_t288 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_1_0_t289 = FSM_dct_8x8_stage_1_0_t288[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t290 = FSM_dct_8x8_stage_1_0_t289 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_1_0_t291 = FSM_dct_8x8_stage_1_0_t290[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t292 = FSM_dct_8x8_stage_1_0_t291[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t293 = FSM_dct_8x8_stage_1_0_t287;
    FSM_dct_8x8_stage_1_0_t293[FSM_dct_8x8_stage_1_0_t292 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t226 - FSM_dct_8x8_stage_1_0_t232;
    FSM_dct_8x8_stage_1_0_t294 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_1_0_t295 = FSM_dct_8x8_stage_1_0_t294[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t296 = FSM_dct_8x8_stage_1_0_t295 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_1_0_t297 = FSM_dct_8x8_stage_1_0_t296[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t298 = FSM_dct_8x8_stage_1_0_t297[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t299 = FSM_dct_8x8_stage_1_0_t293;
    FSM_dct_8x8_stage_1_0_t299[FSM_dct_8x8_stage_1_0_t298 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t206 - FSM_dct_8x8_stage_1_0_t212;
    FSM_dct_8x8_stage_1_0_t300 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_1_0_t301 = FSM_dct_8x8_stage_1_0_t300[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t302 = FSM_dct_8x8_stage_1_0_t301[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t303 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_1_0_t304 = FSM_dct_8x8_stage_1_0_t303[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t305 = FSM_dct_8x8_stage_1_0_t304[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t306 = i_data_in[FSM_dct_8x8_stage_1_0_t305 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t307 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_1_0_t308 = FSM_dct_8x8_stage_1_0_t307[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t309 = FSM_dct_8x8_stage_1_0_t308 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_1_0_t310 = FSM_dct_8x8_stage_1_0_t309[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t311 = FSM_dct_8x8_stage_1_0_t310[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t312 = i_data_in[FSM_dct_8x8_stage_1_0_t311 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t313 = FSM_dct_8x8_stage_1_0_t306 + FSM_dct_8x8_stage_1_0_t312;
    FSM_dct_8x8_stage_1_0_t314 = FSM_dct_8x8_stage_1_0_t313[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t315 = FSM_dct_8x8_stage_1_0_t299;
    FSM_dct_8x8_stage_1_0_t315[FSM_dct_8x8_stage_1_0_t302 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t314;
    FSM_dct_8x8_stage_1_0_t316 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_1_0_t317 = FSM_dct_8x8_stage_1_0_t316[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t318 = FSM_dct_8x8_stage_1_0_t317 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_1_0_t319 = FSM_dct_8x8_stage_1_0_t318[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t320 = FSM_dct_8x8_stage_1_0_t319[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t321 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_1_0_t322 = FSM_dct_8x8_stage_1_0_t321[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t323 = FSM_dct_8x8_stage_1_0_t322 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_1_0_t324 = FSM_dct_8x8_stage_1_0_t323[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t325 = FSM_dct_8x8_stage_1_0_t324[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t326 = i_data_in[FSM_dct_8x8_stage_1_0_t325 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t327 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_1_0_t328 = FSM_dct_8x8_stage_1_0_t327[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t329 = FSM_dct_8x8_stage_1_0_t328 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_1_0_t330 = FSM_dct_8x8_stage_1_0_t329[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t331 = FSM_dct_8x8_stage_1_0_t330[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t332 = i_data_in[FSM_dct_8x8_stage_1_0_t331 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t333 = FSM_dct_8x8_stage_1_0_t326 + FSM_dct_8x8_stage_1_0_t332;
    FSM_dct_8x8_stage_1_0_t334 = FSM_dct_8x8_stage_1_0_t333[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t335 = FSM_dct_8x8_stage_1_0_t315;
    FSM_dct_8x8_stage_1_0_t335[FSM_dct_8x8_stage_1_0_t320 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t334;
    FSM_dct_8x8_stage_1_0_t336 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_1_0_t337 = FSM_dct_8x8_stage_1_0_t336[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t338 = FSM_dct_8x8_stage_1_0_t337 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_1_0_t339 = FSM_dct_8x8_stage_1_0_t338[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t340 = FSM_dct_8x8_stage_1_0_t339[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t341 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_1_0_t342 = FSM_dct_8x8_stage_1_0_t341[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t343 = FSM_dct_8x8_stage_1_0_t342 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_1_0_t344 = FSM_dct_8x8_stage_1_0_t343[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t345 = FSM_dct_8x8_stage_1_0_t344[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t346 = i_data_in[FSM_dct_8x8_stage_1_0_t345 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t347 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_1_0_t348 = FSM_dct_8x8_stage_1_0_t347[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t349 = FSM_dct_8x8_stage_1_0_t348 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_1_0_t350 = FSM_dct_8x8_stage_1_0_t349[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t351 = FSM_dct_8x8_stage_1_0_t350[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t352 = i_data_in[FSM_dct_8x8_stage_1_0_t351 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t353 = FSM_dct_8x8_stage_1_0_t346 + FSM_dct_8x8_stage_1_0_t352;
    FSM_dct_8x8_stage_1_0_t354 = FSM_dct_8x8_stage_1_0_t353[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t355 = FSM_dct_8x8_stage_1_0_t335;
    FSM_dct_8x8_stage_1_0_t355[FSM_dct_8x8_stage_1_0_t340 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t354;
    FSM_dct_8x8_stage_1_0_t356 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_1_0_t357 = FSM_dct_8x8_stage_1_0_t356[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t358 = FSM_dct_8x8_stage_1_0_t357 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_1_0_t359 = FSM_dct_8x8_stage_1_0_t358[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t360 = FSM_dct_8x8_stage_1_0_t359[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t361 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_1_0_t362 = FSM_dct_8x8_stage_1_0_t361[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t363 = FSM_dct_8x8_stage_1_0_t362 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_1_0_t364 = FSM_dct_8x8_stage_1_0_t363[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t365 = FSM_dct_8x8_stage_1_0_t364[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t366 = i_data_in[FSM_dct_8x8_stage_1_0_t365 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t367 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_1_0_t368 = FSM_dct_8x8_stage_1_0_t367[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t369 = FSM_dct_8x8_stage_1_0_t368 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_1_0_t370 = FSM_dct_8x8_stage_1_0_t369[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t371 = FSM_dct_8x8_stage_1_0_t370[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t372 = i_data_in[FSM_dct_8x8_stage_1_0_t371 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t373 = FSM_dct_8x8_stage_1_0_t366 + FSM_dct_8x8_stage_1_0_t372;
    FSM_dct_8x8_stage_1_0_t374 = FSM_dct_8x8_stage_1_0_t373[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t375 = FSM_dct_8x8_stage_1_0_t355;
    FSM_dct_8x8_stage_1_0_t375[FSM_dct_8x8_stage_1_0_t360 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t374;
    FSM_dct_8x8_stage_1_0_t376 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_1_0_t377 = FSM_dct_8x8_stage_1_0_t376[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t378 = FSM_dct_8x8_stage_1_0_t377 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_1_0_t379 = FSM_dct_8x8_stage_1_0_t378[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t380 = FSM_dct_8x8_stage_1_0_t379[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t381 = FSM_dct_8x8_stage_1_0_t375;
    FSM_dct_8x8_stage_1_0_t381[FSM_dct_8x8_stage_1_0_t380 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t366 - FSM_dct_8x8_stage_1_0_t372;
    FSM_dct_8x8_stage_1_0_t382 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_1_0_t383 = FSM_dct_8x8_stage_1_0_t382[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t384 = FSM_dct_8x8_stage_1_0_t383 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_1_0_t385 = FSM_dct_8x8_stage_1_0_t384[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t386 = FSM_dct_8x8_stage_1_0_t385[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t387 = FSM_dct_8x8_stage_1_0_t381;
    FSM_dct_8x8_stage_1_0_t387[FSM_dct_8x8_stage_1_0_t386 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t346 - FSM_dct_8x8_stage_1_0_t352;
    FSM_dct_8x8_stage_1_0_t388 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_1_0_t389 = FSM_dct_8x8_stage_1_0_t388[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t390 = FSM_dct_8x8_stage_1_0_t389 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_1_0_t391 = FSM_dct_8x8_stage_1_0_t390[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t392 = FSM_dct_8x8_stage_1_0_t391[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t393 = FSM_dct_8x8_stage_1_0_t387;
    FSM_dct_8x8_stage_1_0_t393[FSM_dct_8x8_stage_1_0_t392 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t326 - FSM_dct_8x8_stage_1_0_t332;
    FSM_dct_8x8_stage_1_0_t394 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_1_0_t395 = FSM_dct_8x8_stage_1_0_t394[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t396 = FSM_dct_8x8_stage_1_0_t395 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_1_0_t397 = FSM_dct_8x8_stage_1_0_t396[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t398 = FSM_dct_8x8_stage_1_0_t397[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t399 = FSM_dct_8x8_stage_1_0_t393;
    FSM_dct_8x8_stage_1_0_t399[FSM_dct_8x8_stage_1_0_t398 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t306 - FSM_dct_8x8_stage_1_0_t312;
    FSM_dct_8x8_stage_1_0_t400 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_1_0_t401 = FSM_dct_8x8_stage_1_0_t400[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t402 = FSM_dct_8x8_stage_1_0_t401[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t403 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_1_0_t404 = FSM_dct_8x8_stage_1_0_t403[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t405 = FSM_dct_8x8_stage_1_0_t404[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t406 = i_data_in[FSM_dct_8x8_stage_1_0_t405 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t407 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_1_0_t408 = FSM_dct_8x8_stage_1_0_t407[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t409 = FSM_dct_8x8_stage_1_0_t408 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_1_0_t410 = FSM_dct_8x8_stage_1_0_t409[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t411 = FSM_dct_8x8_stage_1_0_t410[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t412 = i_data_in[FSM_dct_8x8_stage_1_0_t411 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t413 = FSM_dct_8x8_stage_1_0_t406 + FSM_dct_8x8_stage_1_0_t412;
    FSM_dct_8x8_stage_1_0_t414 = FSM_dct_8x8_stage_1_0_t413[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t415 = FSM_dct_8x8_stage_1_0_t399;
    FSM_dct_8x8_stage_1_0_t415[FSM_dct_8x8_stage_1_0_t402 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t414;
    FSM_dct_8x8_stage_1_0_t416 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_1_0_t417 = FSM_dct_8x8_stage_1_0_t416[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t418 = FSM_dct_8x8_stage_1_0_t417 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_1_0_t419 = FSM_dct_8x8_stage_1_0_t418[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t420 = FSM_dct_8x8_stage_1_0_t419[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t421 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_1_0_t422 = FSM_dct_8x8_stage_1_0_t421[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t423 = FSM_dct_8x8_stage_1_0_t422 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_1_0_t424 = FSM_dct_8x8_stage_1_0_t423[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t425 = FSM_dct_8x8_stage_1_0_t424[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t426 = i_data_in[FSM_dct_8x8_stage_1_0_t425 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t427 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_1_0_t428 = FSM_dct_8x8_stage_1_0_t427[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t429 = FSM_dct_8x8_stage_1_0_t428 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_1_0_t430 = FSM_dct_8x8_stage_1_0_t429[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t431 = FSM_dct_8x8_stage_1_0_t430[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t432 = i_data_in[FSM_dct_8x8_stage_1_0_t431 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t433 = FSM_dct_8x8_stage_1_0_t426 + FSM_dct_8x8_stage_1_0_t432;
    FSM_dct_8x8_stage_1_0_t434 = FSM_dct_8x8_stage_1_0_t433[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t435 = FSM_dct_8x8_stage_1_0_t415;
    FSM_dct_8x8_stage_1_0_t435[FSM_dct_8x8_stage_1_0_t420 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t434;
    FSM_dct_8x8_stage_1_0_t436 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_1_0_t437 = FSM_dct_8x8_stage_1_0_t436[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t438 = FSM_dct_8x8_stage_1_0_t437 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_1_0_t439 = FSM_dct_8x8_stage_1_0_t438[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t440 = FSM_dct_8x8_stage_1_0_t439[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t441 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_1_0_t442 = FSM_dct_8x8_stage_1_0_t441[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t443 = FSM_dct_8x8_stage_1_0_t442 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_1_0_t444 = FSM_dct_8x8_stage_1_0_t443[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t445 = FSM_dct_8x8_stage_1_0_t444[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t446 = i_data_in[FSM_dct_8x8_stage_1_0_t445 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t447 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_1_0_t448 = FSM_dct_8x8_stage_1_0_t447[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t449 = FSM_dct_8x8_stage_1_0_t448 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_1_0_t450 = FSM_dct_8x8_stage_1_0_t449[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t451 = FSM_dct_8x8_stage_1_0_t450[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t452 = i_data_in[FSM_dct_8x8_stage_1_0_t451 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t453 = FSM_dct_8x8_stage_1_0_t446 + FSM_dct_8x8_stage_1_0_t452;
    FSM_dct_8x8_stage_1_0_t454 = FSM_dct_8x8_stage_1_0_t453[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t455 = FSM_dct_8x8_stage_1_0_t435;
    FSM_dct_8x8_stage_1_0_t455[FSM_dct_8x8_stage_1_0_t440 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t454;
    FSM_dct_8x8_stage_1_0_t456 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_1_0_t457 = FSM_dct_8x8_stage_1_0_t456[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t458 = FSM_dct_8x8_stage_1_0_t457 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_1_0_t459 = FSM_dct_8x8_stage_1_0_t458[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t460 = FSM_dct_8x8_stage_1_0_t459[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t461 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_1_0_t462 = FSM_dct_8x8_stage_1_0_t461[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t463 = FSM_dct_8x8_stage_1_0_t462 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_1_0_t464 = FSM_dct_8x8_stage_1_0_t463[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t465 = FSM_dct_8x8_stage_1_0_t464[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t466 = i_data_in[FSM_dct_8x8_stage_1_0_t465 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t467 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_1_0_t468 = FSM_dct_8x8_stage_1_0_t467[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t469 = FSM_dct_8x8_stage_1_0_t468 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_1_0_t470 = FSM_dct_8x8_stage_1_0_t469[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t471 = FSM_dct_8x8_stage_1_0_t470[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t472 = i_data_in[FSM_dct_8x8_stage_1_0_t471 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t473 = FSM_dct_8x8_stage_1_0_t466 + FSM_dct_8x8_stage_1_0_t472;
    FSM_dct_8x8_stage_1_0_t474 = FSM_dct_8x8_stage_1_0_t473[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t475 = FSM_dct_8x8_stage_1_0_t455;
    FSM_dct_8x8_stage_1_0_t475[FSM_dct_8x8_stage_1_0_t460 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t474;
    FSM_dct_8x8_stage_1_0_t476 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_1_0_t477 = FSM_dct_8x8_stage_1_0_t476[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t478 = FSM_dct_8x8_stage_1_0_t477 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_1_0_t479 = FSM_dct_8x8_stage_1_0_t478[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t480 = FSM_dct_8x8_stage_1_0_t479[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t481 = FSM_dct_8x8_stage_1_0_t475;
    FSM_dct_8x8_stage_1_0_t481[FSM_dct_8x8_stage_1_0_t480 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t466 - FSM_dct_8x8_stage_1_0_t472;
    FSM_dct_8x8_stage_1_0_t482 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_1_0_t483 = FSM_dct_8x8_stage_1_0_t482[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t484 = FSM_dct_8x8_stage_1_0_t483 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_1_0_t485 = FSM_dct_8x8_stage_1_0_t484[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t486 = FSM_dct_8x8_stage_1_0_t485[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t487 = FSM_dct_8x8_stage_1_0_t481;
    FSM_dct_8x8_stage_1_0_t487[FSM_dct_8x8_stage_1_0_t486 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t446 - FSM_dct_8x8_stage_1_0_t452;
    FSM_dct_8x8_stage_1_0_t488 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_1_0_t489 = FSM_dct_8x8_stage_1_0_t488[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t490 = FSM_dct_8x8_stage_1_0_t489 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_1_0_t491 = FSM_dct_8x8_stage_1_0_t490[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t492 = FSM_dct_8x8_stage_1_0_t491[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t493 = FSM_dct_8x8_stage_1_0_t487;
    FSM_dct_8x8_stage_1_0_t493[FSM_dct_8x8_stage_1_0_t492 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t426 - FSM_dct_8x8_stage_1_0_t432;
    FSM_dct_8x8_stage_1_0_t494 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_1_0_t495 = FSM_dct_8x8_stage_1_0_t494[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t496 = FSM_dct_8x8_stage_1_0_t495 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_1_0_t497 = FSM_dct_8x8_stage_1_0_t496[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t498 = FSM_dct_8x8_stage_1_0_t497[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t499 = FSM_dct_8x8_stage_1_0_t493;
    FSM_dct_8x8_stage_1_0_t499[FSM_dct_8x8_stage_1_0_t498 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t406 - FSM_dct_8x8_stage_1_0_t412;
    FSM_dct_8x8_stage_1_0_t500 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_1_0_t501 = FSM_dct_8x8_stage_1_0_t500[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t502 = FSM_dct_8x8_stage_1_0_t501[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t503 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_1_0_t504 = FSM_dct_8x8_stage_1_0_t503[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t505 = FSM_dct_8x8_stage_1_0_t504[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t506 = i_data_in[FSM_dct_8x8_stage_1_0_t505 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t507 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_1_0_t508 = FSM_dct_8x8_stage_1_0_t507[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t509 = FSM_dct_8x8_stage_1_0_t508 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_1_0_t510 = FSM_dct_8x8_stage_1_0_t509[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t511 = FSM_dct_8x8_stage_1_0_t510[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t512 = i_data_in[FSM_dct_8x8_stage_1_0_t511 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t513 = FSM_dct_8x8_stage_1_0_t506 + FSM_dct_8x8_stage_1_0_t512;
    FSM_dct_8x8_stage_1_0_t514 = FSM_dct_8x8_stage_1_0_t513[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t515 = FSM_dct_8x8_stage_1_0_t499;
    FSM_dct_8x8_stage_1_0_t515[FSM_dct_8x8_stage_1_0_t502 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t514;
    FSM_dct_8x8_stage_1_0_t516 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_1_0_t517 = FSM_dct_8x8_stage_1_0_t516[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t518 = FSM_dct_8x8_stage_1_0_t517 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_1_0_t519 = FSM_dct_8x8_stage_1_0_t518[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t520 = FSM_dct_8x8_stage_1_0_t519[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t521 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_1_0_t522 = FSM_dct_8x8_stage_1_0_t521[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t523 = FSM_dct_8x8_stage_1_0_t522 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_1_0_t524 = FSM_dct_8x8_stage_1_0_t523[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t525 = FSM_dct_8x8_stage_1_0_t524[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t526 = i_data_in[FSM_dct_8x8_stage_1_0_t525 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t527 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_1_0_t528 = FSM_dct_8x8_stage_1_0_t527[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t529 = FSM_dct_8x8_stage_1_0_t528 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_1_0_t530 = FSM_dct_8x8_stage_1_0_t529[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t531 = FSM_dct_8x8_stage_1_0_t530[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t532 = i_data_in[FSM_dct_8x8_stage_1_0_t531 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t533 = FSM_dct_8x8_stage_1_0_t526 + FSM_dct_8x8_stage_1_0_t532;
    FSM_dct_8x8_stage_1_0_t534 = FSM_dct_8x8_stage_1_0_t533[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t535 = FSM_dct_8x8_stage_1_0_t515;
    FSM_dct_8x8_stage_1_0_t535[FSM_dct_8x8_stage_1_0_t520 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t534;
    FSM_dct_8x8_stage_1_0_t536 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_1_0_t537 = FSM_dct_8x8_stage_1_0_t536[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t538 = FSM_dct_8x8_stage_1_0_t537 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_1_0_t539 = FSM_dct_8x8_stage_1_0_t538[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t540 = FSM_dct_8x8_stage_1_0_t539[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t541 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_1_0_t542 = FSM_dct_8x8_stage_1_0_t541[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t543 = FSM_dct_8x8_stage_1_0_t542 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_1_0_t544 = FSM_dct_8x8_stage_1_0_t543[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t545 = FSM_dct_8x8_stage_1_0_t544[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t546 = i_data_in[FSM_dct_8x8_stage_1_0_t545 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t547 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_1_0_t548 = FSM_dct_8x8_stage_1_0_t547[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t549 = FSM_dct_8x8_stage_1_0_t548 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_1_0_t550 = FSM_dct_8x8_stage_1_0_t549[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t551 = FSM_dct_8x8_stage_1_0_t550[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t552 = i_data_in[FSM_dct_8x8_stage_1_0_t551 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t553 = FSM_dct_8x8_stage_1_0_t546 + FSM_dct_8x8_stage_1_0_t552;
    FSM_dct_8x8_stage_1_0_t554 = FSM_dct_8x8_stage_1_0_t553[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t555 = FSM_dct_8x8_stage_1_0_t535;
    FSM_dct_8x8_stage_1_0_t555[FSM_dct_8x8_stage_1_0_t540 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t554;
    FSM_dct_8x8_stage_1_0_t556 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_1_0_t557 = FSM_dct_8x8_stage_1_0_t556[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t558 = FSM_dct_8x8_stage_1_0_t557 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_1_0_t559 = FSM_dct_8x8_stage_1_0_t558[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t560 = FSM_dct_8x8_stage_1_0_t559[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t561 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_1_0_t562 = FSM_dct_8x8_stage_1_0_t561[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t563 = FSM_dct_8x8_stage_1_0_t562 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_1_0_t564 = FSM_dct_8x8_stage_1_0_t563[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t565 = FSM_dct_8x8_stage_1_0_t564[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t566 = i_data_in[FSM_dct_8x8_stage_1_0_t565 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t567 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_1_0_t568 = FSM_dct_8x8_stage_1_0_t567[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t569 = FSM_dct_8x8_stage_1_0_t568 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_1_0_t570 = FSM_dct_8x8_stage_1_0_t569[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t571 = FSM_dct_8x8_stage_1_0_t570[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t572 = i_data_in[FSM_dct_8x8_stage_1_0_t571 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t573 = FSM_dct_8x8_stage_1_0_t566 + FSM_dct_8x8_stage_1_0_t572;
    FSM_dct_8x8_stage_1_0_t574 = FSM_dct_8x8_stage_1_0_t573[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t575 = FSM_dct_8x8_stage_1_0_t555;
    FSM_dct_8x8_stage_1_0_t575[FSM_dct_8x8_stage_1_0_t560 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t574;
    FSM_dct_8x8_stage_1_0_t576 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_1_0_t577 = FSM_dct_8x8_stage_1_0_t576[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t578 = FSM_dct_8x8_stage_1_0_t577 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_1_0_t579 = FSM_dct_8x8_stage_1_0_t578[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t580 = FSM_dct_8x8_stage_1_0_t579[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t581 = FSM_dct_8x8_stage_1_0_t575;
    FSM_dct_8x8_stage_1_0_t581[FSM_dct_8x8_stage_1_0_t580 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t566 - FSM_dct_8x8_stage_1_0_t572;
    FSM_dct_8x8_stage_1_0_t582 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_1_0_t583 = FSM_dct_8x8_stage_1_0_t582[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t584 = FSM_dct_8x8_stage_1_0_t583 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_1_0_t585 = FSM_dct_8x8_stage_1_0_t584[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t586 = FSM_dct_8x8_stage_1_0_t585[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t587 = FSM_dct_8x8_stage_1_0_t581;
    FSM_dct_8x8_stage_1_0_t587[FSM_dct_8x8_stage_1_0_t586 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t546 - FSM_dct_8x8_stage_1_0_t552;
    FSM_dct_8x8_stage_1_0_t588 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_1_0_t589 = FSM_dct_8x8_stage_1_0_t588[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t590 = FSM_dct_8x8_stage_1_0_t589 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_1_0_t591 = FSM_dct_8x8_stage_1_0_t590[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t592 = FSM_dct_8x8_stage_1_0_t591[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t593 = FSM_dct_8x8_stage_1_0_t587;
    FSM_dct_8x8_stage_1_0_t593[FSM_dct_8x8_stage_1_0_t592 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t526 - FSM_dct_8x8_stage_1_0_t532;
    FSM_dct_8x8_stage_1_0_t594 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_1_0_t595 = FSM_dct_8x8_stage_1_0_t594[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t596 = FSM_dct_8x8_stage_1_0_t595 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_1_0_t597 = FSM_dct_8x8_stage_1_0_t596[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t598 = FSM_dct_8x8_stage_1_0_t597[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t599 = FSM_dct_8x8_stage_1_0_t593;
    FSM_dct_8x8_stage_1_0_t599[FSM_dct_8x8_stage_1_0_t598 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t506 - FSM_dct_8x8_stage_1_0_t512;
    FSM_dct_8x8_stage_1_0_t600 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_1_0_t601 = FSM_dct_8x8_stage_1_0_t600[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t602 = FSM_dct_8x8_stage_1_0_t601[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t603 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_1_0_t604 = FSM_dct_8x8_stage_1_0_t603[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t605 = FSM_dct_8x8_stage_1_0_t604[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t606 = i_data_in[FSM_dct_8x8_stage_1_0_t605 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t607 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_1_0_t608 = FSM_dct_8x8_stage_1_0_t607[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t609 = FSM_dct_8x8_stage_1_0_t608 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_1_0_t610 = FSM_dct_8x8_stage_1_0_t609[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t611 = FSM_dct_8x8_stage_1_0_t610[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t612 = i_data_in[FSM_dct_8x8_stage_1_0_t611 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t613 = FSM_dct_8x8_stage_1_0_t606 + FSM_dct_8x8_stage_1_0_t612;
    FSM_dct_8x8_stage_1_0_t614 = FSM_dct_8x8_stage_1_0_t613[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t615 = FSM_dct_8x8_stage_1_0_t599;
    FSM_dct_8x8_stage_1_0_t615[FSM_dct_8x8_stage_1_0_t602 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t614;
    FSM_dct_8x8_stage_1_0_t616 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_1_0_t617 = FSM_dct_8x8_stage_1_0_t616[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t618 = FSM_dct_8x8_stage_1_0_t617 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_1_0_t619 = FSM_dct_8x8_stage_1_0_t618[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t620 = FSM_dct_8x8_stage_1_0_t619[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t621 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_1_0_t622 = FSM_dct_8x8_stage_1_0_t621[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t623 = FSM_dct_8x8_stage_1_0_t622 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_1_0_t624 = FSM_dct_8x8_stage_1_0_t623[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t625 = FSM_dct_8x8_stage_1_0_t624[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t626 = i_data_in[FSM_dct_8x8_stage_1_0_t625 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t627 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_1_0_t628 = FSM_dct_8x8_stage_1_0_t627[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t629 = FSM_dct_8x8_stage_1_0_t628 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_1_0_t630 = FSM_dct_8x8_stage_1_0_t629[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t631 = FSM_dct_8x8_stage_1_0_t630[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t632 = i_data_in[FSM_dct_8x8_stage_1_0_t631 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t633 = FSM_dct_8x8_stage_1_0_t626 + FSM_dct_8x8_stage_1_0_t632;
    FSM_dct_8x8_stage_1_0_t634 = FSM_dct_8x8_stage_1_0_t633[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t635 = FSM_dct_8x8_stage_1_0_t615;
    FSM_dct_8x8_stage_1_0_t635[FSM_dct_8x8_stage_1_0_t620 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t634;
    FSM_dct_8x8_stage_1_0_t636 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_1_0_t637 = FSM_dct_8x8_stage_1_0_t636[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t638 = FSM_dct_8x8_stage_1_0_t637 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_1_0_t639 = FSM_dct_8x8_stage_1_0_t638[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t640 = FSM_dct_8x8_stage_1_0_t639[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t641 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_1_0_t642 = FSM_dct_8x8_stage_1_0_t641[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t643 = FSM_dct_8x8_stage_1_0_t642 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_1_0_t644 = FSM_dct_8x8_stage_1_0_t643[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t645 = FSM_dct_8x8_stage_1_0_t644[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t646 = i_data_in[FSM_dct_8x8_stage_1_0_t645 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t647 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_1_0_t648 = FSM_dct_8x8_stage_1_0_t647[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t649 = FSM_dct_8x8_stage_1_0_t648 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_1_0_t650 = FSM_dct_8x8_stage_1_0_t649[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t651 = FSM_dct_8x8_stage_1_0_t650[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t652 = i_data_in[FSM_dct_8x8_stage_1_0_t651 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t653 = FSM_dct_8x8_stage_1_0_t646 + FSM_dct_8x8_stage_1_0_t652;
    FSM_dct_8x8_stage_1_0_t654 = FSM_dct_8x8_stage_1_0_t653[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t655 = FSM_dct_8x8_stage_1_0_t635;
    FSM_dct_8x8_stage_1_0_t655[FSM_dct_8x8_stage_1_0_t640 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t654;
    FSM_dct_8x8_stage_1_0_t656 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_1_0_t657 = FSM_dct_8x8_stage_1_0_t656[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t658 = FSM_dct_8x8_stage_1_0_t657 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_1_0_t659 = FSM_dct_8x8_stage_1_0_t658[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t660 = FSM_dct_8x8_stage_1_0_t659[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t661 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_1_0_t662 = FSM_dct_8x8_stage_1_0_t661[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t663 = FSM_dct_8x8_stage_1_0_t662 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_1_0_t664 = FSM_dct_8x8_stage_1_0_t663[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t665 = FSM_dct_8x8_stage_1_0_t664[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t666 = i_data_in[FSM_dct_8x8_stage_1_0_t665 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t667 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_1_0_t668 = FSM_dct_8x8_stage_1_0_t667[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t669 = FSM_dct_8x8_stage_1_0_t668 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_1_0_t670 = FSM_dct_8x8_stage_1_0_t669[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t671 = FSM_dct_8x8_stage_1_0_t670[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t672 = i_data_in[FSM_dct_8x8_stage_1_0_t671 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t673 = FSM_dct_8x8_stage_1_0_t666 + FSM_dct_8x8_stage_1_0_t672;
    FSM_dct_8x8_stage_1_0_t674 = FSM_dct_8x8_stage_1_0_t673[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t675 = FSM_dct_8x8_stage_1_0_t655;
    FSM_dct_8x8_stage_1_0_t675[FSM_dct_8x8_stage_1_0_t660 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t674;
    FSM_dct_8x8_stage_1_0_t676 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_1_0_t677 = FSM_dct_8x8_stage_1_0_t676[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t678 = FSM_dct_8x8_stage_1_0_t677 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_1_0_t679 = FSM_dct_8x8_stage_1_0_t678[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t680 = FSM_dct_8x8_stage_1_0_t679[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t681 = FSM_dct_8x8_stage_1_0_t675;
    FSM_dct_8x8_stage_1_0_t681[FSM_dct_8x8_stage_1_0_t680 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t666 - FSM_dct_8x8_stage_1_0_t672;
    FSM_dct_8x8_stage_1_0_t682 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_1_0_t683 = FSM_dct_8x8_stage_1_0_t682[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t684 = FSM_dct_8x8_stage_1_0_t683 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_1_0_t685 = FSM_dct_8x8_stage_1_0_t684[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t686 = FSM_dct_8x8_stage_1_0_t685[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t687 = FSM_dct_8x8_stage_1_0_t681;
    FSM_dct_8x8_stage_1_0_t687[FSM_dct_8x8_stage_1_0_t686 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t646 - FSM_dct_8x8_stage_1_0_t652;
    FSM_dct_8x8_stage_1_0_t688 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_1_0_t689 = FSM_dct_8x8_stage_1_0_t688[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t690 = FSM_dct_8x8_stage_1_0_t689 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_1_0_t691 = FSM_dct_8x8_stage_1_0_t690[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t692 = FSM_dct_8x8_stage_1_0_t691[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t693 = FSM_dct_8x8_stage_1_0_t687;
    FSM_dct_8x8_stage_1_0_t693[FSM_dct_8x8_stage_1_0_t692 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t626 - FSM_dct_8x8_stage_1_0_t632;
    FSM_dct_8x8_stage_1_0_t694 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_1_0_t695 = FSM_dct_8x8_stage_1_0_t694[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t696 = FSM_dct_8x8_stage_1_0_t695 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_1_0_t697 = FSM_dct_8x8_stage_1_0_t696[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t698 = FSM_dct_8x8_stage_1_0_t697[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t699 = FSM_dct_8x8_stage_1_0_t693;
    FSM_dct_8x8_stage_1_0_t699[FSM_dct_8x8_stage_1_0_t698 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t606 - FSM_dct_8x8_stage_1_0_t612;
    FSM_dct_8x8_stage_1_0_t700 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_1_0_t701 = FSM_dct_8x8_stage_1_0_t700[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t702 = FSM_dct_8x8_stage_1_0_t701[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t703 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_1_0_t704 = FSM_dct_8x8_stage_1_0_t703[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t705 = FSM_dct_8x8_stage_1_0_t704[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t706 = i_data_in[FSM_dct_8x8_stage_1_0_t705 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t707 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_1_0_t708 = FSM_dct_8x8_stage_1_0_t707[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t709 = FSM_dct_8x8_stage_1_0_t708 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_1_0_t710 = FSM_dct_8x8_stage_1_0_t709[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t711 = FSM_dct_8x8_stage_1_0_t710[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t712 = i_data_in[FSM_dct_8x8_stage_1_0_t711 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t713 = FSM_dct_8x8_stage_1_0_t706 + FSM_dct_8x8_stage_1_0_t712;
    FSM_dct_8x8_stage_1_0_t714 = FSM_dct_8x8_stage_1_0_t713[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t715 = FSM_dct_8x8_stage_1_0_t699;
    FSM_dct_8x8_stage_1_0_t715[FSM_dct_8x8_stage_1_0_t702 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t714;
    FSM_dct_8x8_stage_1_0_t716 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_1_0_t717 = FSM_dct_8x8_stage_1_0_t716[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t718 = FSM_dct_8x8_stage_1_0_t717 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_1_0_t719 = FSM_dct_8x8_stage_1_0_t718[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t720 = FSM_dct_8x8_stage_1_0_t719[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t721 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_1_0_t722 = FSM_dct_8x8_stage_1_0_t721[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t723 = FSM_dct_8x8_stage_1_0_t722 + 32'b00000000000000000000000000000001;
    FSM_dct_8x8_stage_1_0_t724 = FSM_dct_8x8_stage_1_0_t723[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t725 = FSM_dct_8x8_stage_1_0_t724[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t726 = i_data_in[FSM_dct_8x8_stage_1_0_t725 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t727 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_1_0_t728 = FSM_dct_8x8_stage_1_0_t727[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t729 = FSM_dct_8x8_stage_1_0_t728 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_1_0_t730 = FSM_dct_8x8_stage_1_0_t729[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t731 = FSM_dct_8x8_stage_1_0_t730[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t732 = i_data_in[FSM_dct_8x8_stage_1_0_t731 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t733 = FSM_dct_8x8_stage_1_0_t726 + FSM_dct_8x8_stage_1_0_t732;
    FSM_dct_8x8_stage_1_0_t734 = FSM_dct_8x8_stage_1_0_t733[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t735 = FSM_dct_8x8_stage_1_0_t715;
    FSM_dct_8x8_stage_1_0_t735[FSM_dct_8x8_stage_1_0_t720 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t734;
    FSM_dct_8x8_stage_1_0_t736 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_1_0_t737 = FSM_dct_8x8_stage_1_0_t736[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t738 = FSM_dct_8x8_stage_1_0_t737 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_1_0_t739 = FSM_dct_8x8_stage_1_0_t738[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t740 = FSM_dct_8x8_stage_1_0_t739[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t741 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_1_0_t742 = FSM_dct_8x8_stage_1_0_t741[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t743 = FSM_dct_8x8_stage_1_0_t742 + 32'b00000000000000000000000000000010;
    FSM_dct_8x8_stage_1_0_t744 = FSM_dct_8x8_stage_1_0_t743[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t745 = FSM_dct_8x8_stage_1_0_t744[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t746 = i_data_in[FSM_dct_8x8_stage_1_0_t745 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t747 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_1_0_t748 = FSM_dct_8x8_stage_1_0_t747[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t749 = FSM_dct_8x8_stage_1_0_t748 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_1_0_t750 = FSM_dct_8x8_stage_1_0_t749[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t751 = FSM_dct_8x8_stage_1_0_t750[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t752 = i_data_in[FSM_dct_8x8_stage_1_0_t751 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t753 = FSM_dct_8x8_stage_1_0_t746 + FSM_dct_8x8_stage_1_0_t752;
    FSM_dct_8x8_stage_1_0_t754 = FSM_dct_8x8_stage_1_0_t753[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t755 = FSM_dct_8x8_stage_1_0_t735;
    FSM_dct_8x8_stage_1_0_t755[FSM_dct_8x8_stage_1_0_t740 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t754;
    FSM_dct_8x8_stage_1_0_t756 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_1_0_t757 = FSM_dct_8x8_stage_1_0_t756[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t758 = FSM_dct_8x8_stage_1_0_t757 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_1_0_t759 = FSM_dct_8x8_stage_1_0_t758[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t760 = FSM_dct_8x8_stage_1_0_t759[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t761 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_1_0_t762 = FSM_dct_8x8_stage_1_0_t761[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t763 = FSM_dct_8x8_stage_1_0_t762 + 32'b00000000000000000000000000000011;
    FSM_dct_8x8_stage_1_0_t764 = FSM_dct_8x8_stage_1_0_t763[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t765 = FSM_dct_8x8_stage_1_0_t764[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t766 = i_data_in[FSM_dct_8x8_stage_1_0_t765 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t767 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_1_0_t768 = FSM_dct_8x8_stage_1_0_t767[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t769 = FSM_dct_8x8_stage_1_0_t768 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_1_0_t770 = FSM_dct_8x8_stage_1_0_t769[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t771 = FSM_dct_8x8_stage_1_0_t770[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t772 = i_data_in[FSM_dct_8x8_stage_1_0_t771 * 32 +: 32];
    FSM_dct_8x8_stage_1_0_t773 = FSM_dct_8x8_stage_1_0_t766 + FSM_dct_8x8_stage_1_0_t772;
    FSM_dct_8x8_stage_1_0_t774 = FSM_dct_8x8_stage_1_0_t773[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t775 = FSM_dct_8x8_stage_1_0_t755;
    FSM_dct_8x8_stage_1_0_t775[FSM_dct_8x8_stage_1_0_t760 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t774;
    FSM_dct_8x8_stage_1_0_t776 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_1_0_t777 = FSM_dct_8x8_stage_1_0_t776[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t778 = FSM_dct_8x8_stage_1_0_t777 + 32'b00000000000000000000000000000100;
    FSM_dct_8x8_stage_1_0_t779 = FSM_dct_8x8_stage_1_0_t778[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t780 = FSM_dct_8x8_stage_1_0_t779[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t781 = FSM_dct_8x8_stage_1_0_t775;
    FSM_dct_8x8_stage_1_0_t781[FSM_dct_8x8_stage_1_0_t780 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t766 - FSM_dct_8x8_stage_1_0_t772;
    FSM_dct_8x8_stage_1_0_t782 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_1_0_t783 = FSM_dct_8x8_stage_1_0_t782[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t784 = FSM_dct_8x8_stage_1_0_t783 + 32'b00000000000000000000000000000101;
    FSM_dct_8x8_stage_1_0_t785 = FSM_dct_8x8_stage_1_0_t784[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t786 = FSM_dct_8x8_stage_1_0_t785[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t787 = FSM_dct_8x8_stage_1_0_t781;
    FSM_dct_8x8_stage_1_0_t787[FSM_dct_8x8_stage_1_0_t786 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t746 - FSM_dct_8x8_stage_1_0_t752;
    FSM_dct_8x8_stage_1_0_t788 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_1_0_t789 = FSM_dct_8x8_stage_1_0_t788[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t790 = FSM_dct_8x8_stage_1_0_t789 + 32'b00000000000000000000000000000110;
    FSM_dct_8x8_stage_1_0_t791 = FSM_dct_8x8_stage_1_0_t790[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t792 = FSM_dct_8x8_stage_1_0_t791[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t793 = FSM_dct_8x8_stage_1_0_t787;
    FSM_dct_8x8_stage_1_0_t793[FSM_dct_8x8_stage_1_0_t792 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t726 - FSM_dct_8x8_stage_1_0_t732;
    FSM_dct_8x8_stage_1_0_t794 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_1_0_t795 = FSM_dct_8x8_stage_1_0_t794[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t796 = FSM_dct_8x8_stage_1_0_t795 + 32'b00000000000000000000000000000111;
    FSM_dct_8x8_stage_1_0_t797 = FSM_dct_8x8_stage_1_0_t796[6'b0 * 1 +: 32 * 1];
    FSM_dct_8x8_stage_1_0_t798 = FSM_dct_8x8_stage_1_0_t797[5'b0 * 1 +: 6 * 1];
    FSM_dct_8x8_stage_1_0_t799 = FSM_dct_8x8_stage_1_0_t793;
    FSM_dct_8x8_stage_1_0_t799[FSM_dct_8x8_stage_1_0_t798 * 32 +: 32] = FSM_dct_8x8_stage_1_0_t706 - FSM_dct_8x8_stage_1_0_t712;
end

assign FSM_dct_8x8_stage_1_0_in_ready = 1'b1;

always @(posedge clk) begin
    FSM_dct_8x8_stage_1_0_st_dummy_reg <= FSM_dct_8x8_stage_1_0_st_dummy_reg;
    if (rst) begin
        FSM_dct_8x8_stage_1_0_st_dummy_reg <= 32'b0;
    end
end
/* End submodules of dct_8x8_stage_1 */
/* End module dct_8x8_stage_1 */
endgenerate
endmodule
