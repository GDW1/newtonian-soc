package perf_pkg;
	typedef logic [63:0] counter_t;	
endpackage : perf_pkg