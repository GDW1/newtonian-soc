`timescale 1ns / 1ps

module mix_columns_inner
(
    input wire clk,
    input wire rst,
    input wire [64-1:0] i_data_lower,
    input wire [64-1:0] i_data_higher,
    input wire i_valid,
    output wire i_ready,
    output wire [64-1:0] o_data_out_lower,
    output wire [64-1:0] o_data_out_higher,
    output wire o_valid,
    input wire o_ready
);

generate
/*
    Begin module mix_columns
*/
/*
    Wires declared by mix_columns
*/
wire FSM_mix_columns_0_in_ready;
wire [64-1:0] FSM_mix_columns_0_out_data_out_lower;
wire [64-1:0] FSM_mix_columns_0_out_data_out_higher;
wire FSM_mix_columns_0_out_valid;
/* End wires declared by mix_columns */

/*
    Wiring by mix_columns
*/
assign i_ready = FSM_mix_columns_0_in_ready;
assign o_data_out_lower = FSM_mix_columns_0_out_data_out_lower;
assign o_data_out_higher = FSM_mix_columns_0_out_data_out_higher;
assign o_valid = FSM_mix_columns_0_out_valid;
/* End wiring by mix_columns */

/*
    Submodules of mix_columns
*/
reg [64-1:0] FSM_mix_columns_0_st_dummy_reg = 64'b0;

reg [128-1:0] FSM_mix_columns_0_t0;
reg [64-1:0] FSM_mix_columns_0_t1;
reg [64-1:0] FSM_mix_columns_0_t2;
reg [6-1:0] FSM_mix_columns_0_t3;
reg [128-1:0] FSM_mix_columns_0_t4;
reg [64-1:0] FSM_mix_columns_0_t5;
reg [64-1:0] FSM_mix_columns_0_t6;
reg [6-1:0] FSM_mix_columns_0_t7;
reg [64-1:0] FSM_mix_columns_0_t8;
reg [6-1:0] FSM_mix_columns_0_t9;
reg [128-1:0] FSM_mix_columns_0_t10;
reg [64-1:0] FSM_mix_columns_0_t11;
reg [128-1:0] FSM_mix_columns_0_t12;
reg [64-1:0] FSM_mix_columns_0_t13;
reg [64-1:0] FSM_mix_columns_0_t14;
reg [6-1:0] FSM_mix_columns_0_t15;
reg [128-1:0] FSM_mix_columns_0_t16;
reg [64-1:0] FSM_mix_columns_0_t17;
reg [128-1:0] FSM_mix_columns_0_t18;
reg [64-1:0] FSM_mix_columns_0_t19;
reg [64-1:0] FSM_mix_columns_0_t20;
reg [6-1:0] FSM_mix_columns_0_t21;
reg [128-1:0] FSM_mix_columns_0_t22;
reg [64-1:0] FSM_mix_columns_0_t23;
reg [128-1:0] FSM_mix_columns_0_t24;
reg [64-1:0] FSM_mix_columns_0_t25;
reg [64-1:0] FSM_mix_columns_0_t26;
reg [6-1:0] FSM_mix_columns_0_t27;
reg [64-1:0] FSM_mix_columns_0_t28;
reg [6-1:0] FSM_mix_columns_0_t29;
reg [128-1:0] FSM_mix_columns_0_t30;
reg [64-1:0] FSM_mix_columns_0_t31;
reg [64-1:0] FSM_mix_columns_0_t32;
reg [6-1:0] FSM_mix_columns_0_t33;
reg [128-1:0] FSM_mix_columns_0_t34;
reg [64-1:0] FSM_mix_columns_0_t35;
reg [64-1:0] FSM_mix_columns_0_t36;
reg [6-1:0] FSM_mix_columns_0_t37;
reg [64-1:0] FSM_mix_columns_0_t38;
reg [6-1:0] FSM_mix_columns_0_t39;
reg [64-1:0] FSM_mix_columns_0_t40;
reg [6-1:0] FSM_mix_columns_0_t41;
reg [128-1:0] FSM_mix_columns_0_t42;
reg [64-1:0] FSM_mix_columns_0_t43;
reg [128-1:0] FSM_mix_columns_0_t44;
reg [64-1:0] FSM_mix_columns_0_t45;
reg [64-1:0] FSM_mix_columns_0_t46;
reg [6-1:0] FSM_mix_columns_0_t47;
reg [128-1:0] FSM_mix_columns_0_t48;
reg [64-1:0] FSM_mix_columns_0_t49;
reg [128-1:0] FSM_mix_columns_0_t50;
reg [64-1:0] FSM_mix_columns_0_t51;
reg [64-1:0] FSM_mix_columns_0_t52;
reg [6-1:0] FSM_mix_columns_0_t53;
reg [128-1:0] FSM_mix_columns_0_t54;
reg [64-1:0] FSM_mix_columns_0_t55;
reg [128-1:0] FSM_mix_columns_0_t56;
reg [64-1:0] FSM_mix_columns_0_t57;
reg [64-1:0] FSM_mix_columns_0_t58;
reg [6-1:0] FSM_mix_columns_0_t59;
reg [128-1:0] FSM_mix_columns_0_t60;
reg [64-1:0] FSM_mix_columns_0_t61;
reg [64-1:0] FSM_mix_columns_0_t62;
reg [6-1:0] FSM_mix_columns_0_t63;
reg [128-1:0] FSM_mix_columns_0_t64;
reg [64-1:0] FSM_mix_columns_0_t65;
reg [64-1:0] FSM_mix_columns_0_t66;
reg [6-1:0] FSM_mix_columns_0_t67;
reg [64-1:0] FSM_mix_columns_0_t68;
reg [6-1:0] FSM_mix_columns_0_t69;
reg [128-1:0] FSM_mix_columns_0_t70;
reg [64-1:0] FSM_mix_columns_0_t71;
reg [128-1:0] FSM_mix_columns_0_t72;
reg [64-1:0] FSM_mix_columns_0_t73;
reg [64-1:0] FSM_mix_columns_0_t74;
reg [6-1:0] FSM_mix_columns_0_t75;
reg [128-1:0] FSM_mix_columns_0_t76;
reg [64-1:0] FSM_mix_columns_0_t77;
reg [128-1:0] FSM_mix_columns_0_t78;
reg [64-1:0] FSM_mix_columns_0_t79;
reg [64-1:0] FSM_mix_columns_0_t80;
reg [6-1:0] FSM_mix_columns_0_t81;
reg [128-1:0] FSM_mix_columns_0_t82;
reg [64-1:0] FSM_mix_columns_0_t83;
reg [128-1:0] FSM_mix_columns_0_t84;
reg [64-1:0] FSM_mix_columns_0_t85;
reg [64-1:0] FSM_mix_columns_0_t86;
reg [6-1:0] FSM_mix_columns_0_t87;
reg [64-1:0] FSM_mix_columns_0_t88;
reg [6-1:0] FSM_mix_columns_0_t89;
reg [128-1:0] FSM_mix_columns_0_t90;
reg [64-1:0] FSM_mix_columns_0_t91;
reg [64-1:0] FSM_mix_columns_0_t92;
reg [6-1:0] FSM_mix_columns_0_t93;
reg [128-1:0] FSM_mix_columns_0_t94;
reg [64-1:0] FSM_mix_columns_0_t95;
reg [64-1:0] FSM_mix_columns_0_t96;
reg [6-1:0] FSM_mix_columns_0_t97;
reg [64-1:0] FSM_mix_columns_0_t98;
reg [6-1:0] FSM_mix_columns_0_t99;
reg [64-1:0] FSM_mix_columns_0_t100;
reg [6-1:0] FSM_mix_columns_0_t101;
reg [128-1:0] FSM_mix_columns_0_t102;
reg [64-1:0] FSM_mix_columns_0_t103;
reg [128-1:0] FSM_mix_columns_0_t104;
reg [64-1:0] FSM_mix_columns_0_t105;
reg [64-1:0] FSM_mix_columns_0_t106;
reg [6-1:0] FSM_mix_columns_0_t107;
reg [128-1:0] FSM_mix_columns_0_t108;
reg [64-1:0] FSM_mix_columns_0_t109;
reg [128-1:0] FSM_mix_columns_0_t110;
reg [64-1:0] FSM_mix_columns_0_t111;
reg [64-1:0] FSM_mix_columns_0_t112;
reg [6-1:0] FSM_mix_columns_0_t113;
reg [128-1:0] FSM_mix_columns_0_t114;
reg [64-1:0] FSM_mix_columns_0_t115;
reg [128-1:0] FSM_mix_columns_0_t116;
reg [64-1:0] FSM_mix_columns_0_t117;
reg [64-1:0] FSM_mix_columns_0_t118;
reg [6-1:0] FSM_mix_columns_0_t119;

assign FSM_mix_columns_0_out_data_out_lower = (((((((((FSM_mix_columns_0_t1 ^ FSM_mix_columns_0_t5) ^ ((i_data_lower & 64'b0000000000000000000000000000000000000000111111110000000000000000) >> FSM_mix_columns_0_t7)) ^ ((i_data_lower & 64'b0000000000000000000000000000000011111111000000000000000000000000) >> FSM_mix_columns_0_t9)) | (((((i_data_lower & 64'b0000000000000000000000000000000000000000000000000000000011111111) ^ FSM_mix_columns_0_t11) ^ FSM_mix_columns_0_t13) ^ ((i_data_lower & 64'b0000000000000000000000000000000011111111000000000000000000000000) >> FSM_mix_columns_0_t9)) << FSM_mix_columns_0_t15)) | (((((i_data_lower & 64'b0000000000000000000000000000000000000000000000000000000011111111) ^ ((i_data_lower & 64'b0000000000000000000000000000000000000000000000001111111100000000) >> FSM_mix_columns_0_t3)) ^ FSM_mix_columns_0_t17) ^ FSM_mix_columns_0_t19) << FSM_mix_columns_0_t21)) | ((((FSM_mix_columns_0_t23 ^ ((i_data_lower & 64'b0000000000000000000000000000000000000000000000001111111100000000) >> FSM_mix_columns_0_t3)) ^ ((i_data_lower & 64'b0000000000000000000000000000000000000000111111110000000000000000) >> FSM_mix_columns_0_t7)) ^ FSM_mix_columns_0_t25) << FSM_mix_columns_0_t27)) | ((((FSM_mix_columns_0_t31 ^ FSM_mix_columns_0_t35) ^ ((i_data_lower & 64'b0000000011111111000000000000000000000000000000000000000000000000) >> FSM_mix_columns_0_t37)) ^ ((i_data_lower & 64'b1111111100000000000000000000000000000000000000000000000000000000) >> FSM_mix_columns_0_t39)) << FSM_mix_columns_0_t41)) | ((((((i_data_lower & 64'b0000000000000000000000001111111100000000000000000000000000000000) >> FSM_mix_columns_0_t29) ^ FSM_mix_columns_0_t43) ^ FSM_mix_columns_0_t45) ^ ((i_data_lower & 64'b1111111100000000000000000000000000000000000000000000000000000000) >> FSM_mix_columns_0_t39)) << FSM_mix_columns_0_t47)) | ((((((i_data_lower & 64'b0000000000000000000000001111111100000000000000000000000000000000) >> FSM_mix_columns_0_t29) ^ ((i_data_lower & 64'b0000000000000000111111110000000000000000000000000000000000000000) >> FSM_mix_columns_0_t33)) ^ FSM_mix_columns_0_t49) ^ FSM_mix_columns_0_t51) << FSM_mix_columns_0_t53)) | ((((FSM_mix_columns_0_t55 ^ ((i_data_lower & 64'b0000000000000000111111110000000000000000000000000000000000000000) >> FSM_mix_columns_0_t33)) ^ ((i_data_lower & 64'b0000000011111111000000000000000000000000000000000000000000000000) >> FSM_mix_columns_0_t37)) ^ FSM_mix_columns_0_t57) << FSM_mix_columns_0_t59);
assign FSM_mix_columns_0_out_data_out_higher = (((((((((FSM_mix_columns_0_t61 ^ FSM_mix_columns_0_t65) ^ ((i_data_higher & 64'b0000000000000000000000000000000000000000111111110000000000000000) >> FSM_mix_columns_0_t67)) ^ ((i_data_higher & 64'b0000000000000000000000000000000011111111000000000000000000000000) >> FSM_mix_columns_0_t69)) | (((((i_data_higher & 64'b0000000000000000000000000000000000000000000000000000000011111111) ^ FSM_mix_columns_0_t71) ^ FSM_mix_columns_0_t73) ^ ((i_data_higher & 64'b0000000000000000000000000000000011111111000000000000000000000000) >> FSM_mix_columns_0_t69)) << FSM_mix_columns_0_t75)) | (((((i_data_higher & 64'b0000000000000000000000000000000000000000000000000000000011111111) ^ ((i_data_higher & 64'b0000000000000000000000000000000000000000000000001111111100000000) >> FSM_mix_columns_0_t63)) ^ FSM_mix_columns_0_t77) ^ FSM_mix_columns_0_t79) << FSM_mix_columns_0_t81)) | ((((FSM_mix_columns_0_t83 ^ ((i_data_higher & 64'b0000000000000000000000000000000000000000000000001111111100000000) >> FSM_mix_columns_0_t63)) ^ ((i_data_higher & 64'b0000000000000000000000000000000000000000111111110000000000000000) >> FSM_mix_columns_0_t67)) ^ FSM_mix_columns_0_t85) << FSM_mix_columns_0_t87)) | ((((FSM_mix_columns_0_t91 ^ FSM_mix_columns_0_t95) ^ ((i_data_higher & 64'b0000000011111111000000000000000000000000000000000000000000000000) >> FSM_mix_columns_0_t97)) ^ ((i_data_higher & 64'b1111111100000000000000000000000000000000000000000000000000000000) >> FSM_mix_columns_0_t99)) << FSM_mix_columns_0_t101)) | ((((((i_data_higher & 64'b0000000000000000000000001111111100000000000000000000000000000000) >> FSM_mix_columns_0_t89) ^ FSM_mix_columns_0_t103) ^ FSM_mix_columns_0_t105) ^ ((i_data_higher & 64'b1111111100000000000000000000000000000000000000000000000000000000) >> FSM_mix_columns_0_t99)) << FSM_mix_columns_0_t107)) | ((((((i_data_higher & 64'b0000000000000000000000001111111100000000000000000000000000000000) >> FSM_mix_columns_0_t89) ^ ((i_data_higher & 64'b0000000000000000111111110000000000000000000000000000000000000000) >> FSM_mix_columns_0_t93)) ^ FSM_mix_columns_0_t109) ^ FSM_mix_columns_0_t111) << FSM_mix_columns_0_t113)) | ((((FSM_mix_columns_0_t115 ^ ((i_data_higher & 64'b0000000000000000111111110000000000000000000000000000000000000000) >> FSM_mix_columns_0_t93)) ^ ((i_data_higher & 64'b0000000011111111000000000000000000000000000000000000000000000000) >> FSM_mix_columns_0_t97)) ^ FSM_mix_columns_0_t117) << FSM_mix_columns_0_t119);
assign FSM_mix_columns_0_out_valid = 1'b1;

initial begin
    FSM_mix_columns_0_t0 = (i_data_lower & 64'b0000000000000000000000000000000000000000000000000000000011111111) * 64'b0000000000000000000000000000000000000000000000000000000000000010;
    FSM_mix_columns_0_t1 = FSM_mix_columns_0_t0[7'b0 * 1 +: 64 * 1];
    FSM_mix_columns_0_t2 = 64'b0000000000000000000000000000000000000000000000000000000000001000;
    FSM_mix_columns_0_t3 = FSM_mix_columns_0_t2[6'b0 * 1 +: 6 * 1];
    FSM_mix_columns_0_t4 = ((i_data_lower & 64'b0000000000000000000000000000000000000000000000001111111100000000) >> FSM_mix_columns_0_t3) * 64'b0000000000000000000000000000000000000000000000000000000000000011;
    FSM_mix_columns_0_t5 = FSM_mix_columns_0_t4[7'b0 * 1 +: 64 * 1];
    FSM_mix_columns_0_t6 = 64'b0000000000000000000000000000000000000000000000000000000000010000;
    FSM_mix_columns_0_t7 = FSM_mix_columns_0_t6[6'b0 * 1 +: 6 * 1];
    FSM_mix_columns_0_t8 = 64'b0000000000000000000000000000000000000000000000000000000000011000;
    FSM_mix_columns_0_t9 = FSM_mix_columns_0_t8[6'b0 * 1 +: 6 * 1];
    FSM_mix_columns_0_t10 = ((i_data_lower & 64'b0000000000000000000000000000000000000000000000001111111100000000) >> FSM_mix_columns_0_t3) * 64'b0000000000000000000000000000000000000000000000000000000000000010;
    FSM_mix_columns_0_t11 = FSM_mix_columns_0_t10[7'b0 * 1 +: 64 * 1];
    FSM_mix_columns_0_t12 = ((i_data_lower & 64'b0000000000000000000000000000000000000000111111110000000000000000) >> FSM_mix_columns_0_t7) * 64'b0000000000000000000000000000000000000000000000000000000000000011;
    FSM_mix_columns_0_t13 = FSM_mix_columns_0_t12[7'b0 * 1 +: 64 * 1];
    FSM_mix_columns_0_t14 = 64'b0000000000000000000000000000000000000000000000000000000000001000;
    FSM_mix_columns_0_t15 = FSM_mix_columns_0_t14[6'b0 * 1 +: 6 * 1];
    FSM_mix_columns_0_t16 = ((i_data_lower & 64'b0000000000000000000000000000000000000000111111110000000000000000) >> FSM_mix_columns_0_t7) * 64'b0000000000000000000000000000000000000000000000000000000000000010;
    FSM_mix_columns_0_t17 = FSM_mix_columns_0_t16[7'b0 * 1 +: 64 * 1];
    FSM_mix_columns_0_t18 = ((i_data_lower & 64'b0000000000000000000000000000000011111111000000000000000000000000) >> FSM_mix_columns_0_t9) * 64'b0000000000000000000000000000000000000000000000000000000000000011;
    FSM_mix_columns_0_t19 = FSM_mix_columns_0_t18[7'b0 * 1 +: 64 * 1];
    FSM_mix_columns_0_t20 = 64'b0000000000000000000000000000000000000000000000000000000000010000;
    FSM_mix_columns_0_t21 = FSM_mix_columns_0_t20[6'b0 * 1 +: 6 * 1];
    FSM_mix_columns_0_t22 = (i_data_lower & 64'b0000000000000000000000000000000000000000000000000000000011111111) * 64'b0000000000000000000000000000000000000000000000000000000000000011;
    FSM_mix_columns_0_t23 = FSM_mix_columns_0_t22[7'b0 * 1 +: 64 * 1];
    FSM_mix_columns_0_t24 = ((i_data_lower & 64'b0000000000000000000000000000000011111111000000000000000000000000) >> FSM_mix_columns_0_t9) * 64'b0000000000000000000000000000000000000000000000000000000000000010;
    FSM_mix_columns_0_t25 = FSM_mix_columns_0_t24[7'b0 * 1 +: 64 * 1];
    FSM_mix_columns_0_t26 = 64'b0000000000000000000000000000000000000000000000000000000000011000;
    FSM_mix_columns_0_t27 = FSM_mix_columns_0_t26[6'b0 * 1 +: 6 * 1];
    FSM_mix_columns_0_t28 = 64'b0000000000000000000000000000000000000000000000000000000000100000;
    FSM_mix_columns_0_t29 = FSM_mix_columns_0_t28[6'b0 * 1 +: 6 * 1];
    FSM_mix_columns_0_t30 = ((i_data_lower & 64'b0000000000000000000000001111111100000000000000000000000000000000) >> FSM_mix_columns_0_t29) * 64'b0000000000000000000000000000000000000000000000000000000000000010;
    FSM_mix_columns_0_t31 = FSM_mix_columns_0_t30[7'b0 * 1 +: 64 * 1];
    FSM_mix_columns_0_t32 = 64'b0000000000000000000000000000000000000000000000000000000000101000;
    FSM_mix_columns_0_t33 = FSM_mix_columns_0_t32[6'b0 * 1 +: 6 * 1];
    FSM_mix_columns_0_t34 = ((i_data_lower & 64'b0000000000000000111111110000000000000000000000000000000000000000) >> FSM_mix_columns_0_t33) * 64'b0000000000000000000000000000000000000000000000000000000000000011;
    FSM_mix_columns_0_t35 = FSM_mix_columns_0_t34[7'b0 * 1 +: 64 * 1];
    FSM_mix_columns_0_t36 = 64'b0000000000000000000000000000000000000000000000000000000000110000;
    FSM_mix_columns_0_t37 = FSM_mix_columns_0_t36[6'b0 * 1 +: 6 * 1];
    FSM_mix_columns_0_t38 = 64'b0000000000000000000000000000000000000000000000000000000000111000;
    FSM_mix_columns_0_t39 = FSM_mix_columns_0_t38[6'b0 * 1 +: 6 * 1];
    FSM_mix_columns_0_t40 = 64'b0000000000000000000000000000000000000000000000000000000000100000;
    FSM_mix_columns_0_t41 = FSM_mix_columns_0_t40[6'b0 * 1 +: 6 * 1];
    FSM_mix_columns_0_t42 = ((i_data_lower & 64'b0000000000000000111111110000000000000000000000000000000000000000) >> FSM_mix_columns_0_t33) * 64'b0000000000000000000000000000000000000000000000000000000000000010;
    FSM_mix_columns_0_t43 = FSM_mix_columns_0_t42[7'b0 * 1 +: 64 * 1];
    FSM_mix_columns_0_t44 = ((i_data_lower & 64'b0000000011111111000000000000000000000000000000000000000000000000) >> FSM_mix_columns_0_t37) * 64'b0000000000000000000000000000000000000000000000000000000000000011;
    FSM_mix_columns_0_t45 = FSM_mix_columns_0_t44[7'b0 * 1 +: 64 * 1];
    FSM_mix_columns_0_t46 = 64'b0000000000000000000000000000000000000000000000000000000000101000;
    FSM_mix_columns_0_t47 = FSM_mix_columns_0_t46[6'b0 * 1 +: 6 * 1];
    FSM_mix_columns_0_t48 = ((i_data_lower & 64'b0000000011111111000000000000000000000000000000000000000000000000) >> FSM_mix_columns_0_t37) * 64'b0000000000000000000000000000000000000000000000000000000000000010;
    FSM_mix_columns_0_t49 = FSM_mix_columns_0_t48[7'b0 * 1 +: 64 * 1];
    FSM_mix_columns_0_t50 = ((i_data_lower & 64'b1111111100000000000000000000000000000000000000000000000000000000) >> FSM_mix_columns_0_t39) * 64'b0000000000000000000000000000000000000000000000000000000000000011;
    FSM_mix_columns_0_t51 = FSM_mix_columns_0_t50[7'b0 * 1 +: 64 * 1];
    FSM_mix_columns_0_t52 = 64'b0000000000000000000000000000000000000000000000000000000000110000;
    FSM_mix_columns_0_t53 = FSM_mix_columns_0_t52[6'b0 * 1 +: 6 * 1];
    FSM_mix_columns_0_t54 = ((i_data_lower & 64'b0000000000000000000000001111111100000000000000000000000000000000) >> FSM_mix_columns_0_t29) * 64'b0000000000000000000000000000000000000000000000000000000000000011;
    FSM_mix_columns_0_t55 = FSM_mix_columns_0_t54[7'b0 * 1 +: 64 * 1];
    FSM_mix_columns_0_t56 = ((i_data_lower & 64'b1111111100000000000000000000000000000000000000000000000000000000) >> FSM_mix_columns_0_t39) * 64'b0000000000000000000000000000000000000000000000000000000000000010;
    FSM_mix_columns_0_t57 = FSM_mix_columns_0_t56[7'b0 * 1 +: 64 * 1];
    FSM_mix_columns_0_t58 = 64'b0000000000000000000000000000000000000000000000000000000000111000;
    FSM_mix_columns_0_t59 = FSM_mix_columns_0_t58[6'b0 * 1 +: 6 * 1];
    FSM_mix_columns_0_t60 = (i_data_higher & 64'b0000000000000000000000000000000000000000000000000000000011111111) * 64'b0000000000000000000000000000000000000000000000000000000000000010;
    FSM_mix_columns_0_t61 = FSM_mix_columns_0_t60[7'b0 * 1 +: 64 * 1];
    FSM_mix_columns_0_t62 = 64'b0000000000000000000000000000000000000000000000000000000000001000;
    FSM_mix_columns_0_t63 = FSM_mix_columns_0_t62[6'b0 * 1 +: 6 * 1];
    FSM_mix_columns_0_t64 = ((i_data_higher & 64'b0000000000000000000000000000000000000000000000001111111100000000) >> FSM_mix_columns_0_t63) * 64'b0000000000000000000000000000000000000000000000000000000000000011;
    FSM_mix_columns_0_t65 = FSM_mix_columns_0_t64[7'b0 * 1 +: 64 * 1];
    FSM_mix_columns_0_t66 = 64'b0000000000000000000000000000000000000000000000000000000000010000;
    FSM_mix_columns_0_t67 = FSM_mix_columns_0_t66[6'b0 * 1 +: 6 * 1];
    FSM_mix_columns_0_t68 = 64'b0000000000000000000000000000000000000000000000000000000000011000;
    FSM_mix_columns_0_t69 = FSM_mix_columns_0_t68[6'b0 * 1 +: 6 * 1];
    FSM_mix_columns_0_t70 = ((i_data_higher & 64'b0000000000000000000000000000000000000000000000001111111100000000) >> FSM_mix_columns_0_t63) * 64'b0000000000000000000000000000000000000000000000000000000000000010;
    FSM_mix_columns_0_t71 = FSM_mix_columns_0_t70[7'b0 * 1 +: 64 * 1];
    FSM_mix_columns_0_t72 = ((i_data_higher & 64'b0000000000000000000000000000000000000000111111110000000000000000) >> FSM_mix_columns_0_t67) * 64'b0000000000000000000000000000000000000000000000000000000000000011;
    FSM_mix_columns_0_t73 = FSM_mix_columns_0_t72[7'b0 * 1 +: 64 * 1];
    FSM_mix_columns_0_t74 = 64'b0000000000000000000000000000000000000000000000000000000000001000;
    FSM_mix_columns_0_t75 = FSM_mix_columns_0_t74[6'b0 * 1 +: 6 * 1];
    FSM_mix_columns_0_t76 = ((i_data_higher & 64'b0000000000000000000000000000000000000000111111110000000000000000) >> FSM_mix_columns_0_t67) * 64'b0000000000000000000000000000000000000000000000000000000000000010;
    FSM_mix_columns_0_t77 = FSM_mix_columns_0_t76[7'b0 * 1 +: 64 * 1];
    FSM_mix_columns_0_t78 = ((i_data_higher & 64'b0000000000000000000000000000000011111111000000000000000000000000) >> FSM_mix_columns_0_t69) * 64'b0000000000000000000000000000000000000000000000000000000000000011;
    FSM_mix_columns_0_t79 = FSM_mix_columns_0_t78[7'b0 * 1 +: 64 * 1];
    FSM_mix_columns_0_t80 = 64'b0000000000000000000000000000000000000000000000000000000000010000;
    FSM_mix_columns_0_t81 = FSM_mix_columns_0_t80[6'b0 * 1 +: 6 * 1];
    FSM_mix_columns_0_t82 = (i_data_higher & 64'b0000000000000000000000000000000000000000000000000000000011111111) * 64'b0000000000000000000000000000000000000000000000000000000000000011;
    FSM_mix_columns_0_t83 = FSM_mix_columns_0_t82[7'b0 * 1 +: 64 * 1];
    FSM_mix_columns_0_t84 = ((i_data_higher & 64'b0000000000000000000000000000000011111111000000000000000000000000) >> FSM_mix_columns_0_t69) * 64'b0000000000000000000000000000000000000000000000000000000000000010;
    FSM_mix_columns_0_t85 = FSM_mix_columns_0_t84[7'b0 * 1 +: 64 * 1];
    FSM_mix_columns_0_t86 = 64'b0000000000000000000000000000000000000000000000000000000000011000;
    FSM_mix_columns_0_t87 = FSM_mix_columns_0_t86[6'b0 * 1 +: 6 * 1];
    FSM_mix_columns_0_t88 = 64'b0000000000000000000000000000000000000000000000000000000000100000;
    FSM_mix_columns_0_t89 = FSM_mix_columns_0_t88[6'b0 * 1 +: 6 * 1];
    FSM_mix_columns_0_t90 = ((i_data_higher & 64'b0000000000000000000000001111111100000000000000000000000000000000) >> FSM_mix_columns_0_t89) * 64'b0000000000000000000000000000000000000000000000000000000000000010;
    FSM_mix_columns_0_t91 = FSM_mix_columns_0_t90[7'b0 * 1 +: 64 * 1];
    FSM_mix_columns_0_t92 = 64'b0000000000000000000000000000000000000000000000000000000000101000;
    FSM_mix_columns_0_t93 = FSM_mix_columns_0_t92[6'b0 * 1 +: 6 * 1];
    FSM_mix_columns_0_t94 = ((i_data_higher & 64'b0000000000000000111111110000000000000000000000000000000000000000) >> FSM_mix_columns_0_t93) * 64'b0000000000000000000000000000000000000000000000000000000000000011;
    FSM_mix_columns_0_t95 = FSM_mix_columns_0_t94[7'b0 * 1 +: 64 * 1];
    FSM_mix_columns_0_t96 = 64'b0000000000000000000000000000000000000000000000000000000000110000;
    FSM_mix_columns_0_t97 = FSM_mix_columns_0_t96[6'b0 * 1 +: 6 * 1];
    FSM_mix_columns_0_t98 = 64'b0000000000000000000000000000000000000000000000000000000000111000;
    FSM_mix_columns_0_t99 = FSM_mix_columns_0_t98[6'b0 * 1 +: 6 * 1];
    FSM_mix_columns_0_t100 = 64'b0000000000000000000000000000000000000000000000000000000000100000;
    FSM_mix_columns_0_t101 = FSM_mix_columns_0_t100[6'b0 * 1 +: 6 * 1];
    FSM_mix_columns_0_t102 = ((i_data_higher & 64'b0000000000000000111111110000000000000000000000000000000000000000) >> FSM_mix_columns_0_t93) * 64'b0000000000000000000000000000000000000000000000000000000000000010;
    FSM_mix_columns_0_t103 = FSM_mix_columns_0_t102[7'b0 * 1 +: 64 * 1];
    FSM_mix_columns_0_t104 = ((i_data_higher & 64'b0000000011111111000000000000000000000000000000000000000000000000) >> FSM_mix_columns_0_t97) * 64'b0000000000000000000000000000000000000000000000000000000000000011;
    FSM_mix_columns_0_t105 = FSM_mix_columns_0_t104[7'b0 * 1 +: 64 * 1];
    FSM_mix_columns_0_t106 = 64'b0000000000000000000000000000000000000000000000000000000000101000;
    FSM_mix_columns_0_t107 = FSM_mix_columns_0_t106[6'b0 * 1 +: 6 * 1];
    FSM_mix_columns_0_t108 = ((i_data_higher & 64'b0000000011111111000000000000000000000000000000000000000000000000) >> FSM_mix_columns_0_t97) * 64'b0000000000000000000000000000000000000000000000000000000000000010;
    FSM_mix_columns_0_t109 = FSM_mix_columns_0_t108[7'b0 * 1 +: 64 * 1];
    FSM_mix_columns_0_t110 = ((i_data_higher & 64'b1111111100000000000000000000000000000000000000000000000000000000) >> FSM_mix_columns_0_t99) * 64'b0000000000000000000000000000000000000000000000000000000000000011;
    FSM_mix_columns_0_t111 = FSM_mix_columns_0_t110[7'b0 * 1 +: 64 * 1];
    FSM_mix_columns_0_t112 = 64'b0000000000000000000000000000000000000000000000000000000000110000;
    FSM_mix_columns_0_t113 = FSM_mix_columns_0_t112[6'b0 * 1 +: 6 * 1];
    FSM_mix_columns_0_t114 = ((i_data_higher & 64'b0000000000000000000000001111111100000000000000000000000000000000) >> FSM_mix_columns_0_t89) * 64'b0000000000000000000000000000000000000000000000000000000000000011;
    FSM_mix_columns_0_t115 = FSM_mix_columns_0_t114[7'b0 * 1 +: 64 * 1];
    FSM_mix_columns_0_t116 = ((i_data_higher & 64'b1111111100000000000000000000000000000000000000000000000000000000) >> FSM_mix_columns_0_t99) * 64'b0000000000000000000000000000000000000000000000000000000000000010;
    FSM_mix_columns_0_t117 = FSM_mix_columns_0_t116[7'b0 * 1 +: 64 * 1];
    FSM_mix_columns_0_t118 = 64'b0000000000000000000000000000000000000000000000000000000000111000;
    FSM_mix_columns_0_t119 = FSM_mix_columns_0_t118[6'b0 * 1 +: 6 * 1];
end

always @* begin
    FSM_mix_columns_0_t0 = (i_data_lower & 64'b0000000000000000000000000000000000000000000000000000000011111111) * 64'b0000000000000000000000000000000000000000000000000000000000000010;
    FSM_mix_columns_0_t1 = FSM_mix_columns_0_t0[7'b0 * 1 +: 64 * 1];
    FSM_mix_columns_0_t2 = 64'b0000000000000000000000000000000000000000000000000000000000001000;
    FSM_mix_columns_0_t3 = FSM_mix_columns_0_t2[6'b0 * 1 +: 6 * 1];
    FSM_mix_columns_0_t4 = ((i_data_lower & 64'b0000000000000000000000000000000000000000000000001111111100000000) >> FSM_mix_columns_0_t3) * 64'b0000000000000000000000000000000000000000000000000000000000000011;
    FSM_mix_columns_0_t5 = FSM_mix_columns_0_t4[7'b0 * 1 +: 64 * 1];
    FSM_mix_columns_0_t6 = 64'b0000000000000000000000000000000000000000000000000000000000010000;
    FSM_mix_columns_0_t7 = FSM_mix_columns_0_t6[6'b0 * 1 +: 6 * 1];
    FSM_mix_columns_0_t8 = 64'b0000000000000000000000000000000000000000000000000000000000011000;
    FSM_mix_columns_0_t9 = FSM_mix_columns_0_t8[6'b0 * 1 +: 6 * 1];
    FSM_mix_columns_0_t10 = ((i_data_lower & 64'b0000000000000000000000000000000000000000000000001111111100000000) >> FSM_mix_columns_0_t3) * 64'b0000000000000000000000000000000000000000000000000000000000000010;
    FSM_mix_columns_0_t11 = FSM_mix_columns_0_t10[7'b0 * 1 +: 64 * 1];
    FSM_mix_columns_0_t12 = ((i_data_lower & 64'b0000000000000000000000000000000000000000111111110000000000000000) >> FSM_mix_columns_0_t7) * 64'b0000000000000000000000000000000000000000000000000000000000000011;
    FSM_mix_columns_0_t13 = FSM_mix_columns_0_t12[7'b0 * 1 +: 64 * 1];
    FSM_mix_columns_0_t14 = 64'b0000000000000000000000000000000000000000000000000000000000001000;
    FSM_mix_columns_0_t15 = FSM_mix_columns_0_t14[6'b0 * 1 +: 6 * 1];
    FSM_mix_columns_0_t16 = ((i_data_lower & 64'b0000000000000000000000000000000000000000111111110000000000000000) >> FSM_mix_columns_0_t7) * 64'b0000000000000000000000000000000000000000000000000000000000000010;
    FSM_mix_columns_0_t17 = FSM_mix_columns_0_t16[7'b0 * 1 +: 64 * 1];
    FSM_mix_columns_0_t18 = ((i_data_lower & 64'b0000000000000000000000000000000011111111000000000000000000000000) >> FSM_mix_columns_0_t9) * 64'b0000000000000000000000000000000000000000000000000000000000000011;
    FSM_mix_columns_0_t19 = FSM_mix_columns_0_t18[7'b0 * 1 +: 64 * 1];
    FSM_mix_columns_0_t20 = 64'b0000000000000000000000000000000000000000000000000000000000010000;
    FSM_mix_columns_0_t21 = FSM_mix_columns_0_t20[6'b0 * 1 +: 6 * 1];
    FSM_mix_columns_0_t22 = (i_data_lower & 64'b0000000000000000000000000000000000000000000000000000000011111111) * 64'b0000000000000000000000000000000000000000000000000000000000000011;
    FSM_mix_columns_0_t23 = FSM_mix_columns_0_t22[7'b0 * 1 +: 64 * 1];
    FSM_mix_columns_0_t24 = ((i_data_lower & 64'b0000000000000000000000000000000011111111000000000000000000000000) >> FSM_mix_columns_0_t9) * 64'b0000000000000000000000000000000000000000000000000000000000000010;
    FSM_mix_columns_0_t25 = FSM_mix_columns_0_t24[7'b0 * 1 +: 64 * 1];
    FSM_mix_columns_0_t26 = 64'b0000000000000000000000000000000000000000000000000000000000011000;
    FSM_mix_columns_0_t27 = FSM_mix_columns_0_t26[6'b0 * 1 +: 6 * 1];
    FSM_mix_columns_0_t28 = 64'b0000000000000000000000000000000000000000000000000000000000100000;
    FSM_mix_columns_0_t29 = FSM_mix_columns_0_t28[6'b0 * 1 +: 6 * 1];
    FSM_mix_columns_0_t30 = ((i_data_lower & 64'b0000000000000000000000001111111100000000000000000000000000000000) >> FSM_mix_columns_0_t29) * 64'b0000000000000000000000000000000000000000000000000000000000000010;
    FSM_mix_columns_0_t31 = FSM_mix_columns_0_t30[7'b0 * 1 +: 64 * 1];
    FSM_mix_columns_0_t32 = 64'b0000000000000000000000000000000000000000000000000000000000101000;
    FSM_mix_columns_0_t33 = FSM_mix_columns_0_t32[6'b0 * 1 +: 6 * 1];
    FSM_mix_columns_0_t34 = ((i_data_lower & 64'b0000000000000000111111110000000000000000000000000000000000000000) >> FSM_mix_columns_0_t33) * 64'b0000000000000000000000000000000000000000000000000000000000000011;
    FSM_mix_columns_0_t35 = FSM_mix_columns_0_t34[7'b0 * 1 +: 64 * 1];
    FSM_mix_columns_0_t36 = 64'b0000000000000000000000000000000000000000000000000000000000110000;
    FSM_mix_columns_0_t37 = FSM_mix_columns_0_t36[6'b0 * 1 +: 6 * 1];
    FSM_mix_columns_0_t38 = 64'b0000000000000000000000000000000000000000000000000000000000111000;
    FSM_mix_columns_0_t39 = FSM_mix_columns_0_t38[6'b0 * 1 +: 6 * 1];
    FSM_mix_columns_0_t40 = 64'b0000000000000000000000000000000000000000000000000000000000100000;
    FSM_mix_columns_0_t41 = FSM_mix_columns_0_t40[6'b0 * 1 +: 6 * 1];
    FSM_mix_columns_0_t42 = ((i_data_lower & 64'b0000000000000000111111110000000000000000000000000000000000000000) >> FSM_mix_columns_0_t33) * 64'b0000000000000000000000000000000000000000000000000000000000000010;
    FSM_mix_columns_0_t43 = FSM_mix_columns_0_t42[7'b0 * 1 +: 64 * 1];
    FSM_mix_columns_0_t44 = ((i_data_lower & 64'b0000000011111111000000000000000000000000000000000000000000000000) >> FSM_mix_columns_0_t37) * 64'b0000000000000000000000000000000000000000000000000000000000000011;
    FSM_mix_columns_0_t45 = FSM_mix_columns_0_t44[7'b0 * 1 +: 64 * 1];
    FSM_mix_columns_0_t46 = 64'b0000000000000000000000000000000000000000000000000000000000101000;
    FSM_mix_columns_0_t47 = FSM_mix_columns_0_t46[6'b0 * 1 +: 6 * 1];
    FSM_mix_columns_0_t48 = ((i_data_lower & 64'b0000000011111111000000000000000000000000000000000000000000000000) >> FSM_mix_columns_0_t37) * 64'b0000000000000000000000000000000000000000000000000000000000000010;
    FSM_mix_columns_0_t49 = FSM_mix_columns_0_t48[7'b0 * 1 +: 64 * 1];
    FSM_mix_columns_0_t50 = ((i_data_lower & 64'b1111111100000000000000000000000000000000000000000000000000000000) >> FSM_mix_columns_0_t39) * 64'b0000000000000000000000000000000000000000000000000000000000000011;
    FSM_mix_columns_0_t51 = FSM_mix_columns_0_t50[7'b0 * 1 +: 64 * 1];
    FSM_mix_columns_0_t52 = 64'b0000000000000000000000000000000000000000000000000000000000110000;
    FSM_mix_columns_0_t53 = FSM_mix_columns_0_t52[6'b0 * 1 +: 6 * 1];
    FSM_mix_columns_0_t54 = ((i_data_lower & 64'b0000000000000000000000001111111100000000000000000000000000000000) >> FSM_mix_columns_0_t29) * 64'b0000000000000000000000000000000000000000000000000000000000000011;
    FSM_mix_columns_0_t55 = FSM_mix_columns_0_t54[7'b0 * 1 +: 64 * 1];
    FSM_mix_columns_0_t56 = ((i_data_lower & 64'b1111111100000000000000000000000000000000000000000000000000000000) >> FSM_mix_columns_0_t39) * 64'b0000000000000000000000000000000000000000000000000000000000000010;
    FSM_mix_columns_0_t57 = FSM_mix_columns_0_t56[7'b0 * 1 +: 64 * 1];
    FSM_mix_columns_0_t58 = 64'b0000000000000000000000000000000000000000000000000000000000111000;
    FSM_mix_columns_0_t59 = FSM_mix_columns_0_t58[6'b0 * 1 +: 6 * 1];
    FSM_mix_columns_0_t60 = (i_data_higher & 64'b0000000000000000000000000000000000000000000000000000000011111111) * 64'b0000000000000000000000000000000000000000000000000000000000000010;
    FSM_mix_columns_0_t61 = FSM_mix_columns_0_t60[7'b0 * 1 +: 64 * 1];
    FSM_mix_columns_0_t62 = 64'b0000000000000000000000000000000000000000000000000000000000001000;
    FSM_mix_columns_0_t63 = FSM_mix_columns_0_t62[6'b0 * 1 +: 6 * 1];
    FSM_mix_columns_0_t64 = ((i_data_higher & 64'b0000000000000000000000000000000000000000000000001111111100000000) >> FSM_mix_columns_0_t63) * 64'b0000000000000000000000000000000000000000000000000000000000000011;
    FSM_mix_columns_0_t65 = FSM_mix_columns_0_t64[7'b0 * 1 +: 64 * 1];
    FSM_mix_columns_0_t66 = 64'b0000000000000000000000000000000000000000000000000000000000010000;
    FSM_mix_columns_0_t67 = FSM_mix_columns_0_t66[6'b0 * 1 +: 6 * 1];
    FSM_mix_columns_0_t68 = 64'b0000000000000000000000000000000000000000000000000000000000011000;
    FSM_mix_columns_0_t69 = FSM_mix_columns_0_t68[6'b0 * 1 +: 6 * 1];
    FSM_mix_columns_0_t70 = ((i_data_higher & 64'b0000000000000000000000000000000000000000000000001111111100000000) >> FSM_mix_columns_0_t63) * 64'b0000000000000000000000000000000000000000000000000000000000000010;
    FSM_mix_columns_0_t71 = FSM_mix_columns_0_t70[7'b0 * 1 +: 64 * 1];
    FSM_mix_columns_0_t72 = ((i_data_higher & 64'b0000000000000000000000000000000000000000111111110000000000000000) >> FSM_mix_columns_0_t67) * 64'b0000000000000000000000000000000000000000000000000000000000000011;
    FSM_mix_columns_0_t73 = FSM_mix_columns_0_t72[7'b0 * 1 +: 64 * 1];
    FSM_mix_columns_0_t74 = 64'b0000000000000000000000000000000000000000000000000000000000001000;
    FSM_mix_columns_0_t75 = FSM_mix_columns_0_t74[6'b0 * 1 +: 6 * 1];
    FSM_mix_columns_0_t76 = ((i_data_higher & 64'b0000000000000000000000000000000000000000111111110000000000000000) >> FSM_mix_columns_0_t67) * 64'b0000000000000000000000000000000000000000000000000000000000000010;
    FSM_mix_columns_0_t77 = FSM_mix_columns_0_t76[7'b0 * 1 +: 64 * 1];
    FSM_mix_columns_0_t78 = ((i_data_higher & 64'b0000000000000000000000000000000011111111000000000000000000000000) >> FSM_mix_columns_0_t69) * 64'b0000000000000000000000000000000000000000000000000000000000000011;
    FSM_mix_columns_0_t79 = FSM_mix_columns_0_t78[7'b0 * 1 +: 64 * 1];
    FSM_mix_columns_0_t80 = 64'b0000000000000000000000000000000000000000000000000000000000010000;
    FSM_mix_columns_0_t81 = FSM_mix_columns_0_t80[6'b0 * 1 +: 6 * 1];
    FSM_mix_columns_0_t82 = (i_data_higher & 64'b0000000000000000000000000000000000000000000000000000000011111111) * 64'b0000000000000000000000000000000000000000000000000000000000000011;
    FSM_mix_columns_0_t83 = FSM_mix_columns_0_t82[7'b0 * 1 +: 64 * 1];
    FSM_mix_columns_0_t84 = ((i_data_higher & 64'b0000000000000000000000000000000011111111000000000000000000000000) >> FSM_mix_columns_0_t69) * 64'b0000000000000000000000000000000000000000000000000000000000000010;
    FSM_mix_columns_0_t85 = FSM_mix_columns_0_t84[7'b0 * 1 +: 64 * 1];
    FSM_mix_columns_0_t86 = 64'b0000000000000000000000000000000000000000000000000000000000011000;
    FSM_mix_columns_0_t87 = FSM_mix_columns_0_t86[6'b0 * 1 +: 6 * 1];
    FSM_mix_columns_0_t88 = 64'b0000000000000000000000000000000000000000000000000000000000100000;
    FSM_mix_columns_0_t89 = FSM_mix_columns_0_t88[6'b0 * 1 +: 6 * 1];
    FSM_mix_columns_0_t90 = ((i_data_higher & 64'b0000000000000000000000001111111100000000000000000000000000000000) >> FSM_mix_columns_0_t89) * 64'b0000000000000000000000000000000000000000000000000000000000000010;
    FSM_mix_columns_0_t91 = FSM_mix_columns_0_t90[7'b0 * 1 +: 64 * 1];
    FSM_mix_columns_0_t92 = 64'b0000000000000000000000000000000000000000000000000000000000101000;
    FSM_mix_columns_0_t93 = FSM_mix_columns_0_t92[6'b0 * 1 +: 6 * 1];
    FSM_mix_columns_0_t94 = ((i_data_higher & 64'b0000000000000000111111110000000000000000000000000000000000000000) >> FSM_mix_columns_0_t93) * 64'b0000000000000000000000000000000000000000000000000000000000000011;
    FSM_mix_columns_0_t95 = FSM_mix_columns_0_t94[7'b0 * 1 +: 64 * 1];
    FSM_mix_columns_0_t96 = 64'b0000000000000000000000000000000000000000000000000000000000110000;
    FSM_mix_columns_0_t97 = FSM_mix_columns_0_t96[6'b0 * 1 +: 6 * 1];
    FSM_mix_columns_0_t98 = 64'b0000000000000000000000000000000000000000000000000000000000111000;
    FSM_mix_columns_0_t99 = FSM_mix_columns_0_t98[6'b0 * 1 +: 6 * 1];
    FSM_mix_columns_0_t100 = 64'b0000000000000000000000000000000000000000000000000000000000100000;
    FSM_mix_columns_0_t101 = FSM_mix_columns_0_t100[6'b0 * 1 +: 6 * 1];
    FSM_mix_columns_0_t102 = ((i_data_higher & 64'b0000000000000000111111110000000000000000000000000000000000000000) >> FSM_mix_columns_0_t93) * 64'b0000000000000000000000000000000000000000000000000000000000000010;
    FSM_mix_columns_0_t103 = FSM_mix_columns_0_t102[7'b0 * 1 +: 64 * 1];
    FSM_mix_columns_0_t104 = ((i_data_higher & 64'b0000000011111111000000000000000000000000000000000000000000000000) >> FSM_mix_columns_0_t97) * 64'b0000000000000000000000000000000000000000000000000000000000000011;
    FSM_mix_columns_0_t105 = FSM_mix_columns_0_t104[7'b0 * 1 +: 64 * 1];
    FSM_mix_columns_0_t106 = 64'b0000000000000000000000000000000000000000000000000000000000101000;
    FSM_mix_columns_0_t107 = FSM_mix_columns_0_t106[6'b0 * 1 +: 6 * 1];
    FSM_mix_columns_0_t108 = ((i_data_higher & 64'b0000000011111111000000000000000000000000000000000000000000000000) >> FSM_mix_columns_0_t97) * 64'b0000000000000000000000000000000000000000000000000000000000000010;
    FSM_mix_columns_0_t109 = FSM_mix_columns_0_t108[7'b0 * 1 +: 64 * 1];
    FSM_mix_columns_0_t110 = ((i_data_higher & 64'b1111111100000000000000000000000000000000000000000000000000000000) >> FSM_mix_columns_0_t99) * 64'b0000000000000000000000000000000000000000000000000000000000000011;
    FSM_mix_columns_0_t111 = FSM_mix_columns_0_t110[7'b0 * 1 +: 64 * 1];
    FSM_mix_columns_0_t112 = 64'b0000000000000000000000000000000000000000000000000000000000110000;
    FSM_mix_columns_0_t113 = FSM_mix_columns_0_t112[6'b0 * 1 +: 6 * 1];
    FSM_mix_columns_0_t114 = ((i_data_higher & 64'b0000000000000000000000001111111100000000000000000000000000000000) >> FSM_mix_columns_0_t89) * 64'b0000000000000000000000000000000000000000000000000000000000000011;
    FSM_mix_columns_0_t115 = FSM_mix_columns_0_t114[7'b0 * 1 +: 64 * 1];
    FSM_mix_columns_0_t116 = ((i_data_higher & 64'b1111111100000000000000000000000000000000000000000000000000000000) >> FSM_mix_columns_0_t99) * 64'b0000000000000000000000000000000000000000000000000000000000000010;
    FSM_mix_columns_0_t117 = FSM_mix_columns_0_t116[7'b0 * 1 +: 64 * 1];
    FSM_mix_columns_0_t118 = 64'b0000000000000000000000000000000000000000000000000000000000111000;
    FSM_mix_columns_0_t119 = FSM_mix_columns_0_t118[6'b0 * 1 +: 6 * 1];
end

assign FSM_mix_columns_0_in_ready = 1'b1;

always @(posedge clk) begin
    FSM_mix_columns_0_st_dummy_reg <= FSM_mix_columns_0_st_dummy_reg;
    if (rst) begin
        FSM_mix_columns_0_st_dummy_reg <= 64'b0;
    end
end
/* End submodules of mix_columns */
/* End module mix_columns */
endgenerate
endmodule
