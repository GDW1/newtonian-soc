package translator_pkg;

	// verilog type for page number
	typedef logic [`DCP_PADDR-12-1:0] pn_t;


endpackage : translator_pkg