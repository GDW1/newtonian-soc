`timescale 1ns / 1ps

module fft_64_stage_2_inner
(
    input wire clk,
    input wire rst,
    input wire [2048-1:0] i_data_in_real,
    input wire [2048-1:0] i_data_in_imag,
    input wire i_valid,
    output wire i_ready,
    output wire [2048-1:0] o_data_out_real,
    output wire [2048-1:0] o_data_out_imag,
    output wire o_valid,
    input wire o_ready
);

generate
/*
    Begin module fft_64_stage_2
*/
/*
    Wires declared by fft_64_stage_2
*/
wire FSM_fft_64_stage_2_0_in_ready;
wire FSM_fft_64_stage_2_0_out_valid;
/* End wires declared by fft_64_stage_2 */


/*
    Submodules of fft_64_stage_2
*/
reg [32-1:0] FSM_fft_64_stage_2_0_st_dummy_reg = 32'b0;

reg [64-1:0] FSM_fft_64_stage_2_0_t0;
reg [32-1:0] FSM_fft_64_stage_2_0_t1;
reg [6-1:0] FSM_fft_64_stage_2_0_t2;
reg [6-1:0] FSM_fft_64_stage_2_0_t3;
reg [32-1:0] FSM_fft_64_stage_2_0_t4;
reg [33-1:0] FSM_fft_64_stage_2_0_t5;
reg [32-1:0] FSM_fft_64_stage_2_0_t6;
reg [6-1:0] FSM_fft_64_stage_2_0_t7;
reg [32-1:0] FSM_fft_64_stage_2_0_t8;
reg [33-1:0] FSM_fft_64_stage_2_0_t9;
reg [32-1:0] FSM_fft_64_stage_2_0_t10;
reg [2048-1:0] FSM_fft_64_stage_2_0_t11;
reg [33-1:0] FSM_fft_64_stage_2_0_t12;
reg [32-1:0] FSM_fft_64_stage_2_0_t13;
reg [6-1:0] FSM_fft_64_stage_2_0_t14;
reg [2048-1:0] FSM_fft_64_stage_2_0_t15;
reg [33-1:0] FSM_fft_64_stage_2_0_t16;
reg [32-1:0] FSM_fft_64_stage_2_0_t17;
reg [6-1:0] FSM_fft_64_stage_2_0_t18;
reg [33-1:0] FSM_fft_64_stage_2_0_t19;
reg [32-1:0] FSM_fft_64_stage_2_0_t20;
reg [6-1:0] FSM_fft_64_stage_2_0_t21;
reg [32-1:0] FSM_fft_64_stage_2_0_t22;
reg [33-1:0] FSM_fft_64_stage_2_0_t23;
reg [32-1:0] FSM_fft_64_stage_2_0_t24;
reg [6-1:0] FSM_fft_64_stage_2_0_t25;
reg [32-1:0] FSM_fft_64_stage_2_0_t26;
reg [33-1:0] FSM_fft_64_stage_2_0_t27;
reg [32-1:0] FSM_fft_64_stage_2_0_t28;
reg [2048-1:0] FSM_fft_64_stage_2_0_t29;
reg [33-1:0] FSM_fft_64_stage_2_0_t30;
reg [32-1:0] FSM_fft_64_stage_2_0_t31;
reg [6-1:0] FSM_fft_64_stage_2_0_t32;
reg [2048-1:0] FSM_fft_64_stage_2_0_t33;
reg [64-1:0] FSM_fft_64_stage_2_0_t34;
reg [32-1:0] FSM_fft_64_stage_2_0_t35;
reg [6-1:0] FSM_fft_64_stage_2_0_t36;
reg [6-1:0] FSM_fft_64_stage_2_0_t37;
reg [32-1:0] FSM_fft_64_stage_2_0_t38;
reg [33-1:0] FSM_fft_64_stage_2_0_t39;
reg [32-1:0] FSM_fft_64_stage_2_0_t40;
reg [6-1:0] FSM_fft_64_stage_2_0_t41;
reg [32-1:0] FSM_fft_64_stage_2_0_t42;
reg [33-1:0] FSM_fft_64_stage_2_0_t43;
reg [32-1:0] FSM_fft_64_stage_2_0_t44;
reg [2048-1:0] FSM_fft_64_stage_2_0_t45;
reg [33-1:0] FSM_fft_64_stage_2_0_t46;
reg [32-1:0] FSM_fft_64_stage_2_0_t47;
reg [6-1:0] FSM_fft_64_stage_2_0_t48;
reg [2048-1:0] FSM_fft_64_stage_2_0_t49;
reg [33-1:0] FSM_fft_64_stage_2_0_t50;
reg [32-1:0] FSM_fft_64_stage_2_0_t51;
reg [6-1:0] FSM_fft_64_stage_2_0_t52;
reg [33-1:0] FSM_fft_64_stage_2_0_t53;
reg [32-1:0] FSM_fft_64_stage_2_0_t54;
reg [6-1:0] FSM_fft_64_stage_2_0_t55;
reg [32-1:0] FSM_fft_64_stage_2_0_t56;
reg [33-1:0] FSM_fft_64_stage_2_0_t57;
reg [32-1:0] FSM_fft_64_stage_2_0_t58;
reg [6-1:0] FSM_fft_64_stage_2_0_t59;
reg [32-1:0] FSM_fft_64_stage_2_0_t60;
reg [33-1:0] FSM_fft_64_stage_2_0_t61;
reg [32-1:0] FSM_fft_64_stage_2_0_t62;
reg [2048-1:0] FSM_fft_64_stage_2_0_t63;
reg [33-1:0] FSM_fft_64_stage_2_0_t64;
reg [32-1:0] FSM_fft_64_stage_2_0_t65;
reg [6-1:0] FSM_fft_64_stage_2_0_t66;
reg [2048-1:0] FSM_fft_64_stage_2_0_t67;
reg [64-1:0] FSM_fft_64_stage_2_0_t68;
reg [32-1:0] FSM_fft_64_stage_2_0_t69;
reg [6-1:0] FSM_fft_64_stage_2_0_t70;
reg [6-1:0] FSM_fft_64_stage_2_0_t71;
reg [32-1:0] FSM_fft_64_stage_2_0_t72;
reg [33-1:0] FSM_fft_64_stage_2_0_t73;
reg [32-1:0] FSM_fft_64_stage_2_0_t74;
reg [6-1:0] FSM_fft_64_stage_2_0_t75;
reg [32-1:0] FSM_fft_64_stage_2_0_t76;
reg [33-1:0] FSM_fft_64_stage_2_0_t77;
reg [32-1:0] FSM_fft_64_stage_2_0_t78;
reg [2048-1:0] FSM_fft_64_stage_2_0_t79;
reg [33-1:0] FSM_fft_64_stage_2_0_t80;
reg [32-1:0] FSM_fft_64_stage_2_0_t81;
reg [6-1:0] FSM_fft_64_stage_2_0_t82;
reg [2048-1:0] FSM_fft_64_stage_2_0_t83;
reg [33-1:0] FSM_fft_64_stage_2_0_t84;
reg [32-1:0] FSM_fft_64_stage_2_0_t85;
reg [6-1:0] FSM_fft_64_stage_2_0_t86;
reg [33-1:0] FSM_fft_64_stage_2_0_t87;
reg [32-1:0] FSM_fft_64_stage_2_0_t88;
reg [6-1:0] FSM_fft_64_stage_2_0_t89;
reg [32-1:0] FSM_fft_64_stage_2_0_t90;
reg [33-1:0] FSM_fft_64_stage_2_0_t91;
reg [32-1:0] FSM_fft_64_stage_2_0_t92;
reg [6-1:0] FSM_fft_64_stage_2_0_t93;
reg [32-1:0] FSM_fft_64_stage_2_0_t94;
reg [33-1:0] FSM_fft_64_stage_2_0_t95;
reg [32-1:0] FSM_fft_64_stage_2_0_t96;
reg [2048-1:0] FSM_fft_64_stage_2_0_t97;
reg [33-1:0] FSM_fft_64_stage_2_0_t98;
reg [32-1:0] FSM_fft_64_stage_2_0_t99;
reg [6-1:0] FSM_fft_64_stage_2_0_t100;
reg [2048-1:0] FSM_fft_64_stage_2_0_t101;
reg [64-1:0] FSM_fft_64_stage_2_0_t102;
reg [32-1:0] FSM_fft_64_stage_2_0_t103;
reg [6-1:0] FSM_fft_64_stage_2_0_t104;
reg [6-1:0] FSM_fft_64_stage_2_0_t105;
reg [32-1:0] FSM_fft_64_stage_2_0_t106;
reg [33-1:0] FSM_fft_64_stage_2_0_t107;
reg [32-1:0] FSM_fft_64_stage_2_0_t108;
reg [6-1:0] FSM_fft_64_stage_2_0_t109;
reg [32-1:0] FSM_fft_64_stage_2_0_t110;
reg [33-1:0] FSM_fft_64_stage_2_0_t111;
reg [32-1:0] FSM_fft_64_stage_2_0_t112;
reg [2048-1:0] FSM_fft_64_stage_2_0_t113;
reg [33-1:0] FSM_fft_64_stage_2_0_t114;
reg [32-1:0] FSM_fft_64_stage_2_0_t115;
reg [6-1:0] FSM_fft_64_stage_2_0_t116;
reg [2048-1:0] FSM_fft_64_stage_2_0_t117;
reg [33-1:0] FSM_fft_64_stage_2_0_t118;
reg [32-1:0] FSM_fft_64_stage_2_0_t119;
reg [6-1:0] FSM_fft_64_stage_2_0_t120;
reg [33-1:0] FSM_fft_64_stage_2_0_t121;
reg [32-1:0] FSM_fft_64_stage_2_0_t122;
reg [6-1:0] FSM_fft_64_stage_2_0_t123;
reg [32-1:0] FSM_fft_64_stage_2_0_t124;
reg [33-1:0] FSM_fft_64_stage_2_0_t125;
reg [32-1:0] FSM_fft_64_stage_2_0_t126;
reg [6-1:0] FSM_fft_64_stage_2_0_t127;
reg [32-1:0] FSM_fft_64_stage_2_0_t128;
reg [33-1:0] FSM_fft_64_stage_2_0_t129;
reg [32-1:0] FSM_fft_64_stage_2_0_t130;
reg [2048-1:0] FSM_fft_64_stage_2_0_t131;
reg [33-1:0] FSM_fft_64_stage_2_0_t132;
reg [32-1:0] FSM_fft_64_stage_2_0_t133;
reg [6-1:0] FSM_fft_64_stage_2_0_t134;
reg [2048-1:0] FSM_fft_64_stage_2_0_t135;
reg [64-1:0] FSM_fft_64_stage_2_0_t136;
reg [32-1:0] FSM_fft_64_stage_2_0_t137;
reg [6-1:0] FSM_fft_64_stage_2_0_t138;
reg [6-1:0] FSM_fft_64_stage_2_0_t139;
reg [32-1:0] FSM_fft_64_stage_2_0_t140;
reg [33-1:0] FSM_fft_64_stage_2_0_t141;
reg [32-1:0] FSM_fft_64_stage_2_0_t142;
reg [6-1:0] FSM_fft_64_stage_2_0_t143;
reg [32-1:0] FSM_fft_64_stage_2_0_t144;
reg [33-1:0] FSM_fft_64_stage_2_0_t145;
reg [32-1:0] FSM_fft_64_stage_2_0_t146;
reg [2048-1:0] FSM_fft_64_stage_2_0_t147;
reg [33-1:0] FSM_fft_64_stage_2_0_t148;
reg [32-1:0] FSM_fft_64_stage_2_0_t149;
reg [6-1:0] FSM_fft_64_stage_2_0_t150;
reg [2048-1:0] FSM_fft_64_stage_2_0_t151;
reg [33-1:0] FSM_fft_64_stage_2_0_t152;
reg [32-1:0] FSM_fft_64_stage_2_0_t153;
reg [6-1:0] FSM_fft_64_stage_2_0_t154;
reg [33-1:0] FSM_fft_64_stage_2_0_t155;
reg [32-1:0] FSM_fft_64_stage_2_0_t156;
reg [6-1:0] FSM_fft_64_stage_2_0_t157;
reg [32-1:0] FSM_fft_64_stage_2_0_t158;
reg [33-1:0] FSM_fft_64_stage_2_0_t159;
reg [32-1:0] FSM_fft_64_stage_2_0_t160;
reg [6-1:0] FSM_fft_64_stage_2_0_t161;
reg [32-1:0] FSM_fft_64_stage_2_0_t162;
reg [33-1:0] FSM_fft_64_stage_2_0_t163;
reg [32-1:0] FSM_fft_64_stage_2_0_t164;
reg [2048-1:0] FSM_fft_64_stage_2_0_t165;
reg [33-1:0] FSM_fft_64_stage_2_0_t166;
reg [32-1:0] FSM_fft_64_stage_2_0_t167;
reg [6-1:0] FSM_fft_64_stage_2_0_t168;
reg [2048-1:0] FSM_fft_64_stage_2_0_t169;
reg [64-1:0] FSM_fft_64_stage_2_0_t170;
reg [32-1:0] FSM_fft_64_stage_2_0_t171;
reg [6-1:0] FSM_fft_64_stage_2_0_t172;
reg [6-1:0] FSM_fft_64_stage_2_0_t173;
reg [32-1:0] FSM_fft_64_stage_2_0_t174;
reg [33-1:0] FSM_fft_64_stage_2_0_t175;
reg [32-1:0] FSM_fft_64_stage_2_0_t176;
reg [6-1:0] FSM_fft_64_stage_2_0_t177;
reg [32-1:0] FSM_fft_64_stage_2_0_t178;
reg [33-1:0] FSM_fft_64_stage_2_0_t179;
reg [32-1:0] FSM_fft_64_stage_2_0_t180;
reg [2048-1:0] FSM_fft_64_stage_2_0_t181;
reg [33-1:0] FSM_fft_64_stage_2_0_t182;
reg [32-1:0] FSM_fft_64_stage_2_0_t183;
reg [6-1:0] FSM_fft_64_stage_2_0_t184;
reg [2048-1:0] FSM_fft_64_stage_2_0_t185;
reg [33-1:0] FSM_fft_64_stage_2_0_t186;
reg [32-1:0] FSM_fft_64_stage_2_0_t187;
reg [6-1:0] FSM_fft_64_stage_2_0_t188;
reg [33-1:0] FSM_fft_64_stage_2_0_t189;
reg [32-1:0] FSM_fft_64_stage_2_0_t190;
reg [6-1:0] FSM_fft_64_stage_2_0_t191;
reg [32-1:0] FSM_fft_64_stage_2_0_t192;
reg [33-1:0] FSM_fft_64_stage_2_0_t193;
reg [32-1:0] FSM_fft_64_stage_2_0_t194;
reg [6-1:0] FSM_fft_64_stage_2_0_t195;
reg [32-1:0] FSM_fft_64_stage_2_0_t196;
reg [33-1:0] FSM_fft_64_stage_2_0_t197;
reg [32-1:0] FSM_fft_64_stage_2_0_t198;
reg [2048-1:0] FSM_fft_64_stage_2_0_t199;
reg [33-1:0] FSM_fft_64_stage_2_0_t200;
reg [32-1:0] FSM_fft_64_stage_2_0_t201;
reg [6-1:0] FSM_fft_64_stage_2_0_t202;
reg [2048-1:0] FSM_fft_64_stage_2_0_t203;
reg [64-1:0] FSM_fft_64_stage_2_0_t204;
reg [32-1:0] FSM_fft_64_stage_2_0_t205;
reg [6-1:0] FSM_fft_64_stage_2_0_t206;
reg [6-1:0] FSM_fft_64_stage_2_0_t207;
reg [32-1:0] FSM_fft_64_stage_2_0_t208;
reg [33-1:0] FSM_fft_64_stage_2_0_t209;
reg [32-1:0] FSM_fft_64_stage_2_0_t210;
reg [6-1:0] FSM_fft_64_stage_2_0_t211;
reg [32-1:0] FSM_fft_64_stage_2_0_t212;
reg [33-1:0] FSM_fft_64_stage_2_0_t213;
reg [32-1:0] FSM_fft_64_stage_2_0_t214;
reg [2048-1:0] FSM_fft_64_stage_2_0_t215;
reg [33-1:0] FSM_fft_64_stage_2_0_t216;
reg [32-1:0] FSM_fft_64_stage_2_0_t217;
reg [6-1:0] FSM_fft_64_stage_2_0_t218;
reg [2048-1:0] FSM_fft_64_stage_2_0_t219;
reg [33-1:0] FSM_fft_64_stage_2_0_t220;
reg [32-1:0] FSM_fft_64_stage_2_0_t221;
reg [6-1:0] FSM_fft_64_stage_2_0_t222;
reg [33-1:0] FSM_fft_64_stage_2_0_t223;
reg [32-1:0] FSM_fft_64_stage_2_0_t224;
reg [6-1:0] FSM_fft_64_stage_2_0_t225;
reg [32-1:0] FSM_fft_64_stage_2_0_t226;
reg [33-1:0] FSM_fft_64_stage_2_0_t227;
reg [32-1:0] FSM_fft_64_stage_2_0_t228;
reg [6-1:0] FSM_fft_64_stage_2_0_t229;
reg [32-1:0] FSM_fft_64_stage_2_0_t230;
reg [33-1:0] FSM_fft_64_stage_2_0_t231;
reg [32-1:0] FSM_fft_64_stage_2_0_t232;
reg [2048-1:0] FSM_fft_64_stage_2_0_t233;
reg [33-1:0] FSM_fft_64_stage_2_0_t234;
reg [32-1:0] FSM_fft_64_stage_2_0_t235;
reg [6-1:0] FSM_fft_64_stage_2_0_t236;
reg [2048-1:0] FSM_fft_64_stage_2_0_t237;
reg [64-1:0] FSM_fft_64_stage_2_0_t238;
reg [32-1:0] FSM_fft_64_stage_2_0_t239;
reg [6-1:0] FSM_fft_64_stage_2_0_t240;
reg [6-1:0] FSM_fft_64_stage_2_0_t241;
reg [32-1:0] FSM_fft_64_stage_2_0_t242;
reg [33-1:0] FSM_fft_64_stage_2_0_t243;
reg [32-1:0] FSM_fft_64_stage_2_0_t244;
reg [6-1:0] FSM_fft_64_stage_2_0_t245;
reg [32-1:0] FSM_fft_64_stage_2_0_t246;
reg [33-1:0] FSM_fft_64_stage_2_0_t247;
reg [32-1:0] FSM_fft_64_stage_2_0_t248;
reg [2048-1:0] FSM_fft_64_stage_2_0_t249;
reg [33-1:0] FSM_fft_64_stage_2_0_t250;
reg [32-1:0] FSM_fft_64_stage_2_0_t251;
reg [6-1:0] FSM_fft_64_stage_2_0_t252;
reg [2048-1:0] FSM_fft_64_stage_2_0_t253;
reg [33-1:0] FSM_fft_64_stage_2_0_t254;
reg [32-1:0] FSM_fft_64_stage_2_0_t255;
reg [6-1:0] FSM_fft_64_stage_2_0_t256;
reg [33-1:0] FSM_fft_64_stage_2_0_t257;
reg [32-1:0] FSM_fft_64_stage_2_0_t258;
reg [6-1:0] FSM_fft_64_stage_2_0_t259;
reg [32-1:0] FSM_fft_64_stage_2_0_t260;
reg [33-1:0] FSM_fft_64_stage_2_0_t261;
reg [32-1:0] FSM_fft_64_stage_2_0_t262;
reg [6-1:0] FSM_fft_64_stage_2_0_t263;
reg [32-1:0] FSM_fft_64_stage_2_0_t264;
reg [33-1:0] FSM_fft_64_stage_2_0_t265;
reg [32-1:0] FSM_fft_64_stage_2_0_t266;
reg [2048-1:0] FSM_fft_64_stage_2_0_t267;
reg [33-1:0] FSM_fft_64_stage_2_0_t268;
reg [32-1:0] FSM_fft_64_stage_2_0_t269;
reg [6-1:0] FSM_fft_64_stage_2_0_t270;
reg [2048-1:0] FSM_fft_64_stage_2_0_t271;
reg [64-1:0] FSM_fft_64_stage_2_0_t272;
reg [32-1:0] FSM_fft_64_stage_2_0_t273;
reg [6-1:0] FSM_fft_64_stage_2_0_t274;
reg [6-1:0] FSM_fft_64_stage_2_0_t275;
reg [32-1:0] FSM_fft_64_stage_2_0_t276;
reg [33-1:0] FSM_fft_64_stage_2_0_t277;
reg [32-1:0] FSM_fft_64_stage_2_0_t278;
reg [6-1:0] FSM_fft_64_stage_2_0_t279;
reg [32-1:0] FSM_fft_64_stage_2_0_t280;
reg [33-1:0] FSM_fft_64_stage_2_0_t281;
reg [32-1:0] FSM_fft_64_stage_2_0_t282;
reg [2048-1:0] FSM_fft_64_stage_2_0_t283;
reg [33-1:0] FSM_fft_64_stage_2_0_t284;
reg [32-1:0] FSM_fft_64_stage_2_0_t285;
reg [6-1:0] FSM_fft_64_stage_2_0_t286;
reg [2048-1:0] FSM_fft_64_stage_2_0_t287;
reg [33-1:0] FSM_fft_64_stage_2_0_t288;
reg [32-1:0] FSM_fft_64_stage_2_0_t289;
reg [6-1:0] FSM_fft_64_stage_2_0_t290;
reg [33-1:0] FSM_fft_64_stage_2_0_t291;
reg [32-1:0] FSM_fft_64_stage_2_0_t292;
reg [6-1:0] FSM_fft_64_stage_2_0_t293;
reg [32-1:0] FSM_fft_64_stage_2_0_t294;
reg [33-1:0] FSM_fft_64_stage_2_0_t295;
reg [32-1:0] FSM_fft_64_stage_2_0_t296;
reg [6-1:0] FSM_fft_64_stage_2_0_t297;
reg [32-1:0] FSM_fft_64_stage_2_0_t298;
reg [33-1:0] FSM_fft_64_stage_2_0_t299;
reg [32-1:0] FSM_fft_64_stage_2_0_t300;
reg [2048-1:0] FSM_fft_64_stage_2_0_t301;
reg [33-1:0] FSM_fft_64_stage_2_0_t302;
reg [32-1:0] FSM_fft_64_stage_2_0_t303;
reg [6-1:0] FSM_fft_64_stage_2_0_t304;
reg [2048-1:0] FSM_fft_64_stage_2_0_t305;
reg [64-1:0] FSM_fft_64_stage_2_0_t306;
reg [32-1:0] FSM_fft_64_stage_2_0_t307;
reg [6-1:0] FSM_fft_64_stage_2_0_t308;
reg [6-1:0] FSM_fft_64_stage_2_0_t309;
reg [32-1:0] FSM_fft_64_stage_2_0_t310;
reg [33-1:0] FSM_fft_64_stage_2_0_t311;
reg [32-1:0] FSM_fft_64_stage_2_0_t312;
reg [6-1:0] FSM_fft_64_stage_2_0_t313;
reg [32-1:0] FSM_fft_64_stage_2_0_t314;
reg [33-1:0] FSM_fft_64_stage_2_0_t315;
reg [32-1:0] FSM_fft_64_stage_2_0_t316;
reg [2048-1:0] FSM_fft_64_stage_2_0_t317;
reg [33-1:0] FSM_fft_64_stage_2_0_t318;
reg [32-1:0] FSM_fft_64_stage_2_0_t319;
reg [6-1:0] FSM_fft_64_stage_2_0_t320;
reg [2048-1:0] FSM_fft_64_stage_2_0_t321;
reg [33-1:0] FSM_fft_64_stage_2_0_t322;
reg [32-1:0] FSM_fft_64_stage_2_0_t323;
reg [6-1:0] FSM_fft_64_stage_2_0_t324;
reg [33-1:0] FSM_fft_64_stage_2_0_t325;
reg [32-1:0] FSM_fft_64_stage_2_0_t326;
reg [6-1:0] FSM_fft_64_stage_2_0_t327;
reg [32-1:0] FSM_fft_64_stage_2_0_t328;
reg [33-1:0] FSM_fft_64_stage_2_0_t329;
reg [32-1:0] FSM_fft_64_stage_2_0_t330;
reg [6-1:0] FSM_fft_64_stage_2_0_t331;
reg [32-1:0] FSM_fft_64_stage_2_0_t332;
reg [33-1:0] FSM_fft_64_stage_2_0_t333;
reg [32-1:0] FSM_fft_64_stage_2_0_t334;
reg [2048-1:0] FSM_fft_64_stage_2_0_t335;
reg [33-1:0] FSM_fft_64_stage_2_0_t336;
reg [32-1:0] FSM_fft_64_stage_2_0_t337;
reg [6-1:0] FSM_fft_64_stage_2_0_t338;
reg [2048-1:0] FSM_fft_64_stage_2_0_t339;
reg [64-1:0] FSM_fft_64_stage_2_0_t340;
reg [32-1:0] FSM_fft_64_stage_2_0_t341;
reg [6-1:0] FSM_fft_64_stage_2_0_t342;
reg [6-1:0] FSM_fft_64_stage_2_0_t343;
reg [32-1:0] FSM_fft_64_stage_2_0_t344;
reg [33-1:0] FSM_fft_64_stage_2_0_t345;
reg [32-1:0] FSM_fft_64_stage_2_0_t346;
reg [6-1:0] FSM_fft_64_stage_2_0_t347;
reg [32-1:0] FSM_fft_64_stage_2_0_t348;
reg [33-1:0] FSM_fft_64_stage_2_0_t349;
reg [32-1:0] FSM_fft_64_stage_2_0_t350;
reg [2048-1:0] FSM_fft_64_stage_2_0_t351;
reg [33-1:0] FSM_fft_64_stage_2_0_t352;
reg [32-1:0] FSM_fft_64_stage_2_0_t353;
reg [6-1:0] FSM_fft_64_stage_2_0_t354;
reg [2048-1:0] FSM_fft_64_stage_2_0_t355;
reg [33-1:0] FSM_fft_64_stage_2_0_t356;
reg [32-1:0] FSM_fft_64_stage_2_0_t357;
reg [6-1:0] FSM_fft_64_stage_2_0_t358;
reg [33-1:0] FSM_fft_64_stage_2_0_t359;
reg [32-1:0] FSM_fft_64_stage_2_0_t360;
reg [6-1:0] FSM_fft_64_stage_2_0_t361;
reg [32-1:0] FSM_fft_64_stage_2_0_t362;
reg [33-1:0] FSM_fft_64_stage_2_0_t363;
reg [32-1:0] FSM_fft_64_stage_2_0_t364;
reg [6-1:0] FSM_fft_64_stage_2_0_t365;
reg [32-1:0] FSM_fft_64_stage_2_0_t366;
reg [33-1:0] FSM_fft_64_stage_2_0_t367;
reg [32-1:0] FSM_fft_64_stage_2_0_t368;
reg [2048-1:0] FSM_fft_64_stage_2_0_t369;
reg [33-1:0] FSM_fft_64_stage_2_0_t370;
reg [32-1:0] FSM_fft_64_stage_2_0_t371;
reg [6-1:0] FSM_fft_64_stage_2_0_t372;
reg [2048-1:0] FSM_fft_64_stage_2_0_t373;
reg [64-1:0] FSM_fft_64_stage_2_0_t374;
reg [32-1:0] FSM_fft_64_stage_2_0_t375;
reg [6-1:0] FSM_fft_64_stage_2_0_t376;
reg [6-1:0] FSM_fft_64_stage_2_0_t377;
reg [32-1:0] FSM_fft_64_stage_2_0_t378;
reg [33-1:0] FSM_fft_64_stage_2_0_t379;
reg [32-1:0] FSM_fft_64_stage_2_0_t380;
reg [6-1:0] FSM_fft_64_stage_2_0_t381;
reg [32-1:0] FSM_fft_64_stage_2_0_t382;
reg [33-1:0] FSM_fft_64_stage_2_0_t383;
reg [32-1:0] FSM_fft_64_stage_2_0_t384;
reg [2048-1:0] FSM_fft_64_stage_2_0_t385;
reg [33-1:0] FSM_fft_64_stage_2_0_t386;
reg [32-1:0] FSM_fft_64_stage_2_0_t387;
reg [6-1:0] FSM_fft_64_stage_2_0_t388;
reg [2048-1:0] FSM_fft_64_stage_2_0_t389;
reg [33-1:0] FSM_fft_64_stage_2_0_t390;
reg [32-1:0] FSM_fft_64_stage_2_0_t391;
reg [6-1:0] FSM_fft_64_stage_2_0_t392;
reg [33-1:0] FSM_fft_64_stage_2_0_t393;
reg [32-1:0] FSM_fft_64_stage_2_0_t394;
reg [6-1:0] FSM_fft_64_stage_2_0_t395;
reg [32-1:0] FSM_fft_64_stage_2_0_t396;
reg [33-1:0] FSM_fft_64_stage_2_0_t397;
reg [32-1:0] FSM_fft_64_stage_2_0_t398;
reg [6-1:0] FSM_fft_64_stage_2_0_t399;
reg [32-1:0] FSM_fft_64_stage_2_0_t400;
reg [33-1:0] FSM_fft_64_stage_2_0_t401;
reg [32-1:0] FSM_fft_64_stage_2_0_t402;
reg [2048-1:0] FSM_fft_64_stage_2_0_t403;
reg [33-1:0] FSM_fft_64_stage_2_0_t404;
reg [32-1:0] FSM_fft_64_stage_2_0_t405;
reg [6-1:0] FSM_fft_64_stage_2_0_t406;
reg [2048-1:0] FSM_fft_64_stage_2_0_t407;
reg [64-1:0] FSM_fft_64_stage_2_0_t408;
reg [32-1:0] FSM_fft_64_stage_2_0_t409;
reg [6-1:0] FSM_fft_64_stage_2_0_t410;
reg [6-1:0] FSM_fft_64_stage_2_0_t411;
reg [32-1:0] FSM_fft_64_stage_2_0_t412;
reg [33-1:0] FSM_fft_64_stage_2_0_t413;
reg [32-1:0] FSM_fft_64_stage_2_0_t414;
reg [6-1:0] FSM_fft_64_stage_2_0_t415;
reg [32-1:0] FSM_fft_64_stage_2_0_t416;
reg [33-1:0] FSM_fft_64_stage_2_0_t417;
reg [32-1:0] FSM_fft_64_stage_2_0_t418;
reg [2048-1:0] FSM_fft_64_stage_2_0_t419;
reg [33-1:0] FSM_fft_64_stage_2_0_t420;
reg [32-1:0] FSM_fft_64_stage_2_0_t421;
reg [6-1:0] FSM_fft_64_stage_2_0_t422;
reg [2048-1:0] FSM_fft_64_stage_2_0_t423;
reg [33-1:0] FSM_fft_64_stage_2_0_t424;
reg [32-1:0] FSM_fft_64_stage_2_0_t425;
reg [6-1:0] FSM_fft_64_stage_2_0_t426;
reg [33-1:0] FSM_fft_64_stage_2_0_t427;
reg [32-1:0] FSM_fft_64_stage_2_0_t428;
reg [6-1:0] FSM_fft_64_stage_2_0_t429;
reg [32-1:0] FSM_fft_64_stage_2_0_t430;
reg [33-1:0] FSM_fft_64_stage_2_0_t431;
reg [32-1:0] FSM_fft_64_stage_2_0_t432;
reg [6-1:0] FSM_fft_64_stage_2_0_t433;
reg [32-1:0] FSM_fft_64_stage_2_0_t434;
reg [33-1:0] FSM_fft_64_stage_2_0_t435;
reg [32-1:0] FSM_fft_64_stage_2_0_t436;
reg [2048-1:0] FSM_fft_64_stage_2_0_t437;
reg [33-1:0] FSM_fft_64_stage_2_0_t438;
reg [32-1:0] FSM_fft_64_stage_2_0_t439;
reg [6-1:0] FSM_fft_64_stage_2_0_t440;
reg [2048-1:0] FSM_fft_64_stage_2_0_t441;
reg [64-1:0] FSM_fft_64_stage_2_0_t442;
reg [32-1:0] FSM_fft_64_stage_2_0_t443;
reg [6-1:0] FSM_fft_64_stage_2_0_t444;
reg [6-1:0] FSM_fft_64_stage_2_0_t445;
reg [32-1:0] FSM_fft_64_stage_2_0_t446;
reg [33-1:0] FSM_fft_64_stage_2_0_t447;
reg [32-1:0] FSM_fft_64_stage_2_0_t448;
reg [6-1:0] FSM_fft_64_stage_2_0_t449;
reg [32-1:0] FSM_fft_64_stage_2_0_t450;
reg [33-1:0] FSM_fft_64_stage_2_0_t451;
reg [32-1:0] FSM_fft_64_stage_2_0_t452;
reg [2048-1:0] FSM_fft_64_stage_2_0_t453;
reg [33-1:0] FSM_fft_64_stage_2_0_t454;
reg [32-1:0] FSM_fft_64_stage_2_0_t455;
reg [6-1:0] FSM_fft_64_stage_2_0_t456;
reg [2048-1:0] FSM_fft_64_stage_2_0_t457;
reg [33-1:0] FSM_fft_64_stage_2_0_t458;
reg [32-1:0] FSM_fft_64_stage_2_0_t459;
reg [6-1:0] FSM_fft_64_stage_2_0_t460;
reg [33-1:0] FSM_fft_64_stage_2_0_t461;
reg [32-1:0] FSM_fft_64_stage_2_0_t462;
reg [6-1:0] FSM_fft_64_stage_2_0_t463;
reg [32-1:0] FSM_fft_64_stage_2_0_t464;
reg [33-1:0] FSM_fft_64_stage_2_0_t465;
reg [32-1:0] FSM_fft_64_stage_2_0_t466;
reg [6-1:0] FSM_fft_64_stage_2_0_t467;
reg [32-1:0] FSM_fft_64_stage_2_0_t468;
reg [33-1:0] FSM_fft_64_stage_2_0_t469;
reg [32-1:0] FSM_fft_64_stage_2_0_t470;
reg [2048-1:0] FSM_fft_64_stage_2_0_t471;
reg [33-1:0] FSM_fft_64_stage_2_0_t472;
reg [32-1:0] FSM_fft_64_stage_2_0_t473;
reg [6-1:0] FSM_fft_64_stage_2_0_t474;
reg [2048-1:0] FSM_fft_64_stage_2_0_t475;
reg [64-1:0] FSM_fft_64_stage_2_0_t476;
reg [32-1:0] FSM_fft_64_stage_2_0_t477;
reg [6-1:0] FSM_fft_64_stage_2_0_t478;
reg [6-1:0] FSM_fft_64_stage_2_0_t479;
reg [32-1:0] FSM_fft_64_stage_2_0_t480;
reg [33-1:0] FSM_fft_64_stage_2_0_t481;
reg [32-1:0] FSM_fft_64_stage_2_0_t482;
reg [6-1:0] FSM_fft_64_stage_2_0_t483;
reg [32-1:0] FSM_fft_64_stage_2_0_t484;
reg [33-1:0] FSM_fft_64_stage_2_0_t485;
reg [32-1:0] FSM_fft_64_stage_2_0_t486;
reg [2048-1:0] FSM_fft_64_stage_2_0_t487;
reg [33-1:0] FSM_fft_64_stage_2_0_t488;
reg [32-1:0] FSM_fft_64_stage_2_0_t489;
reg [6-1:0] FSM_fft_64_stage_2_0_t490;
reg [2048-1:0] FSM_fft_64_stage_2_0_t491;
reg [33-1:0] FSM_fft_64_stage_2_0_t492;
reg [32-1:0] FSM_fft_64_stage_2_0_t493;
reg [6-1:0] FSM_fft_64_stage_2_0_t494;
reg [33-1:0] FSM_fft_64_stage_2_0_t495;
reg [32-1:0] FSM_fft_64_stage_2_0_t496;
reg [6-1:0] FSM_fft_64_stage_2_0_t497;
reg [32-1:0] FSM_fft_64_stage_2_0_t498;
reg [33-1:0] FSM_fft_64_stage_2_0_t499;
reg [32-1:0] FSM_fft_64_stage_2_0_t500;
reg [6-1:0] FSM_fft_64_stage_2_0_t501;
reg [32-1:0] FSM_fft_64_stage_2_0_t502;
reg [33-1:0] FSM_fft_64_stage_2_0_t503;
reg [32-1:0] FSM_fft_64_stage_2_0_t504;
reg [2048-1:0] FSM_fft_64_stage_2_0_t505;
reg [33-1:0] FSM_fft_64_stage_2_0_t506;
reg [32-1:0] FSM_fft_64_stage_2_0_t507;
reg [6-1:0] FSM_fft_64_stage_2_0_t508;
reg [2048-1:0] FSM_fft_64_stage_2_0_t509;
reg [64-1:0] FSM_fft_64_stage_2_0_t510;
reg [32-1:0] FSM_fft_64_stage_2_0_t511;
reg [6-1:0] FSM_fft_64_stage_2_0_t512;
reg [6-1:0] FSM_fft_64_stage_2_0_t513;
reg [32-1:0] FSM_fft_64_stage_2_0_t514;
reg [33-1:0] FSM_fft_64_stage_2_0_t515;
reg [32-1:0] FSM_fft_64_stage_2_0_t516;
reg [6-1:0] FSM_fft_64_stage_2_0_t517;
reg [32-1:0] FSM_fft_64_stage_2_0_t518;
reg [33-1:0] FSM_fft_64_stage_2_0_t519;
reg [32-1:0] FSM_fft_64_stage_2_0_t520;
reg [2048-1:0] FSM_fft_64_stage_2_0_t521;
reg [33-1:0] FSM_fft_64_stage_2_0_t522;
reg [32-1:0] FSM_fft_64_stage_2_0_t523;
reg [6-1:0] FSM_fft_64_stage_2_0_t524;
reg [2048-1:0] FSM_fft_64_stage_2_0_t525;
reg [33-1:0] FSM_fft_64_stage_2_0_t526;
reg [32-1:0] FSM_fft_64_stage_2_0_t527;
reg [6-1:0] FSM_fft_64_stage_2_0_t528;
reg [33-1:0] FSM_fft_64_stage_2_0_t529;
reg [32-1:0] FSM_fft_64_stage_2_0_t530;
reg [6-1:0] FSM_fft_64_stage_2_0_t531;
reg [32-1:0] FSM_fft_64_stage_2_0_t532;
reg [33-1:0] FSM_fft_64_stage_2_0_t533;
reg [32-1:0] FSM_fft_64_stage_2_0_t534;
reg [6-1:0] FSM_fft_64_stage_2_0_t535;
reg [32-1:0] FSM_fft_64_stage_2_0_t536;
reg [33-1:0] FSM_fft_64_stage_2_0_t537;
reg [32-1:0] FSM_fft_64_stage_2_0_t538;
reg [2048-1:0] FSM_fft_64_stage_2_0_t539;
reg [33-1:0] FSM_fft_64_stage_2_0_t540;
reg [32-1:0] FSM_fft_64_stage_2_0_t541;
reg [6-1:0] FSM_fft_64_stage_2_0_t542;
reg [2048-1:0] FSM_fft_64_stage_2_0_t543;
reg [6-1:0] FSM_fft_64_stage_2_0_t544;
reg [6-1:0] FSM_fft_64_stage_2_0_t545;
reg [32-1:0] FSM_fft_64_stage_2_0_t546;
reg [33-1:0] FSM_fft_64_stage_2_0_t547;
reg [32-1:0] FSM_fft_64_stage_2_0_t548;
reg [6-1:0] FSM_fft_64_stage_2_0_t549;
reg [32-1:0] FSM_fft_64_stage_2_0_t550;
reg [33-1:0] FSM_fft_64_stage_2_0_t551;
reg [32-1:0] FSM_fft_64_stage_2_0_t552;
reg [2048-1:0] FSM_fft_64_stage_2_0_t553;
reg [33-1:0] FSM_fft_64_stage_2_0_t554;
reg [32-1:0] FSM_fft_64_stage_2_0_t555;
reg [6-1:0] FSM_fft_64_stage_2_0_t556;
reg [2048-1:0] FSM_fft_64_stage_2_0_t557;
reg [33-1:0] FSM_fft_64_stage_2_0_t558;
reg [32-1:0] FSM_fft_64_stage_2_0_t559;
reg [6-1:0] FSM_fft_64_stage_2_0_t560;
reg [33-1:0] FSM_fft_64_stage_2_0_t561;
reg [32-1:0] FSM_fft_64_stage_2_0_t562;
reg [6-1:0] FSM_fft_64_stage_2_0_t563;
reg [32-1:0] FSM_fft_64_stage_2_0_t564;
reg [33-1:0] FSM_fft_64_stage_2_0_t565;
reg [32-1:0] FSM_fft_64_stage_2_0_t566;
reg [6-1:0] FSM_fft_64_stage_2_0_t567;
reg [32-1:0] FSM_fft_64_stage_2_0_t568;
reg [33-1:0] FSM_fft_64_stage_2_0_t569;
reg [32-1:0] FSM_fft_64_stage_2_0_t570;
reg [2048-1:0] FSM_fft_64_stage_2_0_t571;
reg [33-1:0] FSM_fft_64_stage_2_0_t572;
reg [32-1:0] FSM_fft_64_stage_2_0_t573;
reg [6-1:0] FSM_fft_64_stage_2_0_t574;
reg [2048-1:0] FSM_fft_64_stage_2_0_t575;
reg [6-1:0] FSM_fft_64_stage_2_0_t576;
reg [6-1:0] FSM_fft_64_stage_2_0_t577;
reg [32-1:0] FSM_fft_64_stage_2_0_t578;
reg [33-1:0] FSM_fft_64_stage_2_0_t579;
reg [32-1:0] FSM_fft_64_stage_2_0_t580;
reg [6-1:0] FSM_fft_64_stage_2_0_t581;
reg [32-1:0] FSM_fft_64_stage_2_0_t582;
reg [33-1:0] FSM_fft_64_stage_2_0_t583;
reg [32-1:0] FSM_fft_64_stage_2_0_t584;
reg [2048-1:0] FSM_fft_64_stage_2_0_t585;
reg [33-1:0] FSM_fft_64_stage_2_0_t586;
reg [32-1:0] FSM_fft_64_stage_2_0_t587;
reg [6-1:0] FSM_fft_64_stage_2_0_t588;
reg [2048-1:0] FSM_fft_64_stage_2_0_t589;
reg [33-1:0] FSM_fft_64_stage_2_0_t590;
reg [32-1:0] FSM_fft_64_stage_2_0_t591;
reg [6-1:0] FSM_fft_64_stage_2_0_t592;
reg [33-1:0] FSM_fft_64_stage_2_0_t593;
reg [32-1:0] FSM_fft_64_stage_2_0_t594;
reg [6-1:0] FSM_fft_64_stage_2_0_t595;
reg [32-1:0] FSM_fft_64_stage_2_0_t596;
reg [33-1:0] FSM_fft_64_stage_2_0_t597;
reg [32-1:0] FSM_fft_64_stage_2_0_t598;
reg [6-1:0] FSM_fft_64_stage_2_0_t599;
reg [32-1:0] FSM_fft_64_stage_2_0_t600;
reg [33-1:0] FSM_fft_64_stage_2_0_t601;
reg [32-1:0] FSM_fft_64_stage_2_0_t602;
reg [2048-1:0] FSM_fft_64_stage_2_0_t603;
reg [33-1:0] FSM_fft_64_stage_2_0_t604;
reg [32-1:0] FSM_fft_64_stage_2_0_t605;
reg [6-1:0] FSM_fft_64_stage_2_0_t606;
reg [2048-1:0] FSM_fft_64_stage_2_0_t607;
reg [6-1:0] FSM_fft_64_stage_2_0_t608;
reg [6-1:0] FSM_fft_64_stage_2_0_t609;
reg [32-1:0] FSM_fft_64_stage_2_0_t610;
reg [33-1:0] FSM_fft_64_stage_2_0_t611;
reg [32-1:0] FSM_fft_64_stage_2_0_t612;
reg [6-1:0] FSM_fft_64_stage_2_0_t613;
reg [32-1:0] FSM_fft_64_stage_2_0_t614;
reg [33-1:0] FSM_fft_64_stage_2_0_t615;
reg [32-1:0] FSM_fft_64_stage_2_0_t616;
reg [2048-1:0] FSM_fft_64_stage_2_0_t617;
reg [33-1:0] FSM_fft_64_stage_2_0_t618;
reg [32-1:0] FSM_fft_64_stage_2_0_t619;
reg [6-1:0] FSM_fft_64_stage_2_0_t620;
reg [2048-1:0] FSM_fft_64_stage_2_0_t621;
reg [33-1:0] FSM_fft_64_stage_2_0_t622;
reg [32-1:0] FSM_fft_64_stage_2_0_t623;
reg [6-1:0] FSM_fft_64_stage_2_0_t624;
reg [33-1:0] FSM_fft_64_stage_2_0_t625;
reg [32-1:0] FSM_fft_64_stage_2_0_t626;
reg [6-1:0] FSM_fft_64_stage_2_0_t627;
reg [32-1:0] FSM_fft_64_stage_2_0_t628;
reg [33-1:0] FSM_fft_64_stage_2_0_t629;
reg [32-1:0] FSM_fft_64_stage_2_0_t630;
reg [6-1:0] FSM_fft_64_stage_2_0_t631;
reg [32-1:0] FSM_fft_64_stage_2_0_t632;
reg [33-1:0] FSM_fft_64_stage_2_0_t633;
reg [32-1:0] FSM_fft_64_stage_2_0_t634;
reg [2048-1:0] FSM_fft_64_stage_2_0_t635;
reg [33-1:0] FSM_fft_64_stage_2_0_t636;
reg [32-1:0] FSM_fft_64_stage_2_0_t637;
reg [6-1:0] FSM_fft_64_stage_2_0_t638;
reg [2048-1:0] FSM_fft_64_stage_2_0_t639;
reg [6-1:0] FSM_fft_64_stage_2_0_t640;
reg [6-1:0] FSM_fft_64_stage_2_0_t641;
reg [32-1:0] FSM_fft_64_stage_2_0_t642;
reg [33-1:0] FSM_fft_64_stage_2_0_t643;
reg [32-1:0] FSM_fft_64_stage_2_0_t644;
reg [6-1:0] FSM_fft_64_stage_2_0_t645;
reg [32-1:0] FSM_fft_64_stage_2_0_t646;
reg [33-1:0] FSM_fft_64_stage_2_0_t647;
reg [32-1:0] FSM_fft_64_stage_2_0_t648;
reg [2048-1:0] FSM_fft_64_stage_2_0_t649;
reg [33-1:0] FSM_fft_64_stage_2_0_t650;
reg [32-1:0] FSM_fft_64_stage_2_0_t651;
reg [6-1:0] FSM_fft_64_stage_2_0_t652;
reg [2048-1:0] FSM_fft_64_stage_2_0_t653;
reg [33-1:0] FSM_fft_64_stage_2_0_t654;
reg [32-1:0] FSM_fft_64_stage_2_0_t655;
reg [6-1:0] FSM_fft_64_stage_2_0_t656;
reg [33-1:0] FSM_fft_64_stage_2_0_t657;
reg [32-1:0] FSM_fft_64_stage_2_0_t658;
reg [6-1:0] FSM_fft_64_stage_2_0_t659;
reg [32-1:0] FSM_fft_64_stage_2_0_t660;
reg [33-1:0] FSM_fft_64_stage_2_0_t661;
reg [32-1:0] FSM_fft_64_stage_2_0_t662;
reg [6-1:0] FSM_fft_64_stage_2_0_t663;
reg [32-1:0] FSM_fft_64_stage_2_0_t664;
reg [33-1:0] FSM_fft_64_stage_2_0_t665;
reg [32-1:0] FSM_fft_64_stage_2_0_t666;
reg [2048-1:0] FSM_fft_64_stage_2_0_t667;
reg [33-1:0] FSM_fft_64_stage_2_0_t668;
reg [32-1:0] FSM_fft_64_stage_2_0_t669;
reg [6-1:0] FSM_fft_64_stage_2_0_t670;
reg [2048-1:0] FSM_fft_64_stage_2_0_t671;
reg [6-1:0] FSM_fft_64_stage_2_0_t672;
reg [6-1:0] FSM_fft_64_stage_2_0_t673;
reg [32-1:0] FSM_fft_64_stage_2_0_t674;
reg [33-1:0] FSM_fft_64_stage_2_0_t675;
reg [32-1:0] FSM_fft_64_stage_2_0_t676;
reg [6-1:0] FSM_fft_64_stage_2_0_t677;
reg [32-1:0] FSM_fft_64_stage_2_0_t678;
reg [33-1:0] FSM_fft_64_stage_2_0_t679;
reg [32-1:0] FSM_fft_64_stage_2_0_t680;
reg [2048-1:0] FSM_fft_64_stage_2_0_t681;
reg [33-1:0] FSM_fft_64_stage_2_0_t682;
reg [32-1:0] FSM_fft_64_stage_2_0_t683;
reg [6-1:0] FSM_fft_64_stage_2_0_t684;
reg [2048-1:0] FSM_fft_64_stage_2_0_t685;
reg [33-1:0] FSM_fft_64_stage_2_0_t686;
reg [32-1:0] FSM_fft_64_stage_2_0_t687;
reg [6-1:0] FSM_fft_64_stage_2_0_t688;
reg [33-1:0] FSM_fft_64_stage_2_0_t689;
reg [32-1:0] FSM_fft_64_stage_2_0_t690;
reg [6-1:0] FSM_fft_64_stage_2_0_t691;
reg [32-1:0] FSM_fft_64_stage_2_0_t692;
reg [33-1:0] FSM_fft_64_stage_2_0_t693;
reg [32-1:0] FSM_fft_64_stage_2_0_t694;
reg [6-1:0] FSM_fft_64_stage_2_0_t695;
reg [32-1:0] FSM_fft_64_stage_2_0_t696;
reg [33-1:0] FSM_fft_64_stage_2_0_t697;
reg [32-1:0] FSM_fft_64_stage_2_0_t698;
reg [2048-1:0] FSM_fft_64_stage_2_0_t699;
reg [33-1:0] FSM_fft_64_stage_2_0_t700;
reg [32-1:0] FSM_fft_64_stage_2_0_t701;
reg [6-1:0] FSM_fft_64_stage_2_0_t702;
reg [2048-1:0] FSM_fft_64_stage_2_0_t703;
reg [6-1:0] FSM_fft_64_stage_2_0_t704;
reg [6-1:0] FSM_fft_64_stage_2_0_t705;
reg [32-1:0] FSM_fft_64_stage_2_0_t706;
reg [33-1:0] FSM_fft_64_stage_2_0_t707;
reg [32-1:0] FSM_fft_64_stage_2_0_t708;
reg [6-1:0] FSM_fft_64_stage_2_0_t709;
reg [32-1:0] FSM_fft_64_stage_2_0_t710;
reg [33-1:0] FSM_fft_64_stage_2_0_t711;
reg [32-1:0] FSM_fft_64_stage_2_0_t712;
reg [2048-1:0] FSM_fft_64_stage_2_0_t713;
reg [33-1:0] FSM_fft_64_stage_2_0_t714;
reg [32-1:0] FSM_fft_64_stage_2_0_t715;
reg [6-1:0] FSM_fft_64_stage_2_0_t716;
reg [2048-1:0] FSM_fft_64_stage_2_0_t717;
reg [33-1:0] FSM_fft_64_stage_2_0_t718;
reg [32-1:0] FSM_fft_64_stage_2_0_t719;
reg [6-1:0] FSM_fft_64_stage_2_0_t720;
reg [33-1:0] FSM_fft_64_stage_2_0_t721;
reg [32-1:0] FSM_fft_64_stage_2_0_t722;
reg [6-1:0] FSM_fft_64_stage_2_0_t723;
reg [32-1:0] FSM_fft_64_stage_2_0_t724;
reg [33-1:0] FSM_fft_64_stage_2_0_t725;
reg [32-1:0] FSM_fft_64_stage_2_0_t726;
reg [6-1:0] FSM_fft_64_stage_2_0_t727;
reg [32-1:0] FSM_fft_64_stage_2_0_t728;
reg [33-1:0] FSM_fft_64_stage_2_0_t729;
reg [32-1:0] FSM_fft_64_stage_2_0_t730;
reg [2048-1:0] FSM_fft_64_stage_2_0_t731;
reg [33-1:0] FSM_fft_64_stage_2_0_t732;
reg [32-1:0] FSM_fft_64_stage_2_0_t733;
reg [6-1:0] FSM_fft_64_stage_2_0_t734;
reg [2048-1:0] FSM_fft_64_stage_2_0_t735;
reg [6-1:0] FSM_fft_64_stage_2_0_t736;
reg [6-1:0] FSM_fft_64_stage_2_0_t737;
reg [32-1:0] FSM_fft_64_stage_2_0_t738;
reg [33-1:0] FSM_fft_64_stage_2_0_t739;
reg [32-1:0] FSM_fft_64_stage_2_0_t740;
reg [6-1:0] FSM_fft_64_stage_2_0_t741;
reg [32-1:0] FSM_fft_64_stage_2_0_t742;
reg [33-1:0] FSM_fft_64_stage_2_0_t743;
reg [32-1:0] FSM_fft_64_stage_2_0_t744;
reg [2048-1:0] FSM_fft_64_stage_2_0_t745;
reg [33-1:0] FSM_fft_64_stage_2_0_t746;
reg [32-1:0] FSM_fft_64_stage_2_0_t747;
reg [6-1:0] FSM_fft_64_stage_2_0_t748;
reg [2048-1:0] FSM_fft_64_stage_2_0_t749;
reg [33-1:0] FSM_fft_64_stage_2_0_t750;
reg [32-1:0] FSM_fft_64_stage_2_0_t751;
reg [6-1:0] FSM_fft_64_stage_2_0_t752;
reg [33-1:0] FSM_fft_64_stage_2_0_t753;
reg [32-1:0] FSM_fft_64_stage_2_0_t754;
reg [6-1:0] FSM_fft_64_stage_2_0_t755;
reg [32-1:0] FSM_fft_64_stage_2_0_t756;
reg [33-1:0] FSM_fft_64_stage_2_0_t757;
reg [32-1:0] FSM_fft_64_stage_2_0_t758;
reg [6-1:0] FSM_fft_64_stage_2_0_t759;
reg [32-1:0] FSM_fft_64_stage_2_0_t760;
reg [33-1:0] FSM_fft_64_stage_2_0_t761;
reg [32-1:0] FSM_fft_64_stage_2_0_t762;
reg [2048-1:0] FSM_fft_64_stage_2_0_t763;
reg [33-1:0] FSM_fft_64_stage_2_0_t764;
reg [32-1:0] FSM_fft_64_stage_2_0_t765;
reg [6-1:0] FSM_fft_64_stage_2_0_t766;
reg [2048-1:0] FSM_fft_64_stage_2_0_t767;
reg [6-1:0] FSM_fft_64_stage_2_0_t768;
reg [6-1:0] FSM_fft_64_stage_2_0_t769;
reg [32-1:0] FSM_fft_64_stage_2_0_t770;
reg [33-1:0] FSM_fft_64_stage_2_0_t771;
reg [32-1:0] FSM_fft_64_stage_2_0_t772;
reg [6-1:0] FSM_fft_64_stage_2_0_t773;
reg [32-1:0] FSM_fft_64_stage_2_0_t774;
reg [33-1:0] FSM_fft_64_stage_2_0_t775;
reg [32-1:0] FSM_fft_64_stage_2_0_t776;
reg [2048-1:0] FSM_fft_64_stage_2_0_t777;
reg [33-1:0] FSM_fft_64_stage_2_0_t778;
reg [32-1:0] FSM_fft_64_stage_2_0_t779;
reg [6-1:0] FSM_fft_64_stage_2_0_t780;
reg [2048-1:0] FSM_fft_64_stage_2_0_t781;
reg [33-1:0] FSM_fft_64_stage_2_0_t782;
reg [32-1:0] FSM_fft_64_stage_2_0_t783;
reg [6-1:0] FSM_fft_64_stage_2_0_t784;
reg [33-1:0] FSM_fft_64_stage_2_0_t785;
reg [32-1:0] FSM_fft_64_stage_2_0_t786;
reg [6-1:0] FSM_fft_64_stage_2_0_t787;
reg [32-1:0] FSM_fft_64_stage_2_0_t788;
reg [33-1:0] FSM_fft_64_stage_2_0_t789;
reg [32-1:0] FSM_fft_64_stage_2_0_t790;
reg [6-1:0] FSM_fft_64_stage_2_0_t791;
reg [32-1:0] FSM_fft_64_stage_2_0_t792;
reg [33-1:0] FSM_fft_64_stage_2_0_t793;
reg [32-1:0] FSM_fft_64_stage_2_0_t794;
reg [2048-1:0] FSM_fft_64_stage_2_0_t795;
reg [33-1:0] FSM_fft_64_stage_2_0_t796;
reg [32-1:0] FSM_fft_64_stage_2_0_t797;
reg [6-1:0] FSM_fft_64_stage_2_0_t798;
reg [2048-1:0] FSM_fft_64_stage_2_0_t799;
reg [6-1:0] FSM_fft_64_stage_2_0_t800;
reg [6-1:0] FSM_fft_64_stage_2_0_t801;
reg [32-1:0] FSM_fft_64_stage_2_0_t802;
reg [33-1:0] FSM_fft_64_stage_2_0_t803;
reg [32-1:0] FSM_fft_64_stage_2_0_t804;
reg [6-1:0] FSM_fft_64_stage_2_0_t805;
reg [32-1:0] FSM_fft_64_stage_2_0_t806;
reg [33-1:0] FSM_fft_64_stage_2_0_t807;
reg [32-1:0] FSM_fft_64_stage_2_0_t808;
reg [2048-1:0] FSM_fft_64_stage_2_0_t809;
reg [33-1:0] FSM_fft_64_stage_2_0_t810;
reg [32-1:0] FSM_fft_64_stage_2_0_t811;
reg [6-1:0] FSM_fft_64_stage_2_0_t812;
reg [2048-1:0] FSM_fft_64_stage_2_0_t813;
reg [33-1:0] FSM_fft_64_stage_2_0_t814;
reg [32-1:0] FSM_fft_64_stage_2_0_t815;
reg [6-1:0] FSM_fft_64_stage_2_0_t816;
reg [33-1:0] FSM_fft_64_stage_2_0_t817;
reg [32-1:0] FSM_fft_64_stage_2_0_t818;
reg [6-1:0] FSM_fft_64_stage_2_0_t819;
reg [32-1:0] FSM_fft_64_stage_2_0_t820;
reg [33-1:0] FSM_fft_64_stage_2_0_t821;
reg [32-1:0] FSM_fft_64_stage_2_0_t822;
reg [6-1:0] FSM_fft_64_stage_2_0_t823;
reg [32-1:0] FSM_fft_64_stage_2_0_t824;
reg [33-1:0] FSM_fft_64_stage_2_0_t825;
reg [32-1:0] FSM_fft_64_stage_2_0_t826;
reg [2048-1:0] FSM_fft_64_stage_2_0_t827;
reg [33-1:0] FSM_fft_64_stage_2_0_t828;
reg [32-1:0] FSM_fft_64_stage_2_0_t829;
reg [6-1:0] FSM_fft_64_stage_2_0_t830;
reg [2048-1:0] FSM_fft_64_stage_2_0_t831;
reg [6-1:0] FSM_fft_64_stage_2_0_t832;
reg [6-1:0] FSM_fft_64_stage_2_0_t833;
reg [32-1:0] FSM_fft_64_stage_2_0_t834;
reg [33-1:0] FSM_fft_64_stage_2_0_t835;
reg [32-1:0] FSM_fft_64_stage_2_0_t836;
reg [6-1:0] FSM_fft_64_stage_2_0_t837;
reg [32-1:0] FSM_fft_64_stage_2_0_t838;
reg [33-1:0] FSM_fft_64_stage_2_0_t839;
reg [32-1:0] FSM_fft_64_stage_2_0_t840;
reg [2048-1:0] FSM_fft_64_stage_2_0_t841;
reg [33-1:0] FSM_fft_64_stage_2_0_t842;
reg [32-1:0] FSM_fft_64_stage_2_0_t843;
reg [6-1:0] FSM_fft_64_stage_2_0_t844;
reg [2048-1:0] FSM_fft_64_stage_2_0_t845;
reg [33-1:0] FSM_fft_64_stage_2_0_t846;
reg [32-1:0] FSM_fft_64_stage_2_0_t847;
reg [6-1:0] FSM_fft_64_stage_2_0_t848;
reg [33-1:0] FSM_fft_64_stage_2_0_t849;
reg [32-1:0] FSM_fft_64_stage_2_0_t850;
reg [6-1:0] FSM_fft_64_stage_2_0_t851;
reg [32-1:0] FSM_fft_64_stage_2_0_t852;
reg [33-1:0] FSM_fft_64_stage_2_0_t853;
reg [32-1:0] FSM_fft_64_stage_2_0_t854;
reg [6-1:0] FSM_fft_64_stage_2_0_t855;
reg [32-1:0] FSM_fft_64_stage_2_0_t856;
reg [33-1:0] FSM_fft_64_stage_2_0_t857;
reg [32-1:0] FSM_fft_64_stage_2_0_t858;
reg [2048-1:0] FSM_fft_64_stage_2_0_t859;
reg [33-1:0] FSM_fft_64_stage_2_0_t860;
reg [32-1:0] FSM_fft_64_stage_2_0_t861;
reg [6-1:0] FSM_fft_64_stage_2_0_t862;
reg [2048-1:0] FSM_fft_64_stage_2_0_t863;
reg [6-1:0] FSM_fft_64_stage_2_0_t864;
reg [6-1:0] FSM_fft_64_stage_2_0_t865;
reg [32-1:0] FSM_fft_64_stage_2_0_t866;
reg [33-1:0] FSM_fft_64_stage_2_0_t867;
reg [32-1:0] FSM_fft_64_stage_2_0_t868;
reg [6-1:0] FSM_fft_64_stage_2_0_t869;
reg [32-1:0] FSM_fft_64_stage_2_0_t870;
reg [33-1:0] FSM_fft_64_stage_2_0_t871;
reg [32-1:0] FSM_fft_64_stage_2_0_t872;
reg [2048-1:0] FSM_fft_64_stage_2_0_t873;
reg [33-1:0] FSM_fft_64_stage_2_0_t874;
reg [32-1:0] FSM_fft_64_stage_2_0_t875;
reg [6-1:0] FSM_fft_64_stage_2_0_t876;
reg [2048-1:0] FSM_fft_64_stage_2_0_t877;
reg [33-1:0] FSM_fft_64_stage_2_0_t878;
reg [32-1:0] FSM_fft_64_stage_2_0_t879;
reg [6-1:0] FSM_fft_64_stage_2_0_t880;
reg [33-1:0] FSM_fft_64_stage_2_0_t881;
reg [32-1:0] FSM_fft_64_stage_2_0_t882;
reg [6-1:0] FSM_fft_64_stage_2_0_t883;
reg [32-1:0] FSM_fft_64_stage_2_0_t884;
reg [33-1:0] FSM_fft_64_stage_2_0_t885;
reg [32-1:0] FSM_fft_64_stage_2_0_t886;
reg [6-1:0] FSM_fft_64_stage_2_0_t887;
reg [32-1:0] FSM_fft_64_stage_2_0_t888;
reg [33-1:0] FSM_fft_64_stage_2_0_t889;
reg [32-1:0] FSM_fft_64_stage_2_0_t890;
reg [2048-1:0] FSM_fft_64_stage_2_0_t891;
reg [33-1:0] FSM_fft_64_stage_2_0_t892;
reg [32-1:0] FSM_fft_64_stage_2_0_t893;
reg [6-1:0] FSM_fft_64_stage_2_0_t894;
reg [2048-1:0] FSM_fft_64_stage_2_0_t895;
reg [6-1:0] FSM_fft_64_stage_2_0_t896;
reg [6-1:0] FSM_fft_64_stage_2_0_t897;
reg [32-1:0] FSM_fft_64_stage_2_0_t898;
reg [33-1:0] FSM_fft_64_stage_2_0_t899;
reg [32-1:0] FSM_fft_64_stage_2_0_t900;
reg [6-1:0] FSM_fft_64_stage_2_0_t901;
reg [32-1:0] FSM_fft_64_stage_2_0_t902;
reg [33-1:0] FSM_fft_64_stage_2_0_t903;
reg [32-1:0] FSM_fft_64_stage_2_0_t904;
reg [2048-1:0] FSM_fft_64_stage_2_0_t905;
reg [33-1:0] FSM_fft_64_stage_2_0_t906;
reg [32-1:0] FSM_fft_64_stage_2_0_t907;
reg [6-1:0] FSM_fft_64_stage_2_0_t908;
reg [2048-1:0] FSM_fft_64_stage_2_0_t909;
reg [33-1:0] FSM_fft_64_stage_2_0_t910;
reg [32-1:0] FSM_fft_64_stage_2_0_t911;
reg [6-1:0] FSM_fft_64_stage_2_0_t912;
reg [33-1:0] FSM_fft_64_stage_2_0_t913;
reg [32-1:0] FSM_fft_64_stage_2_0_t914;
reg [6-1:0] FSM_fft_64_stage_2_0_t915;
reg [32-1:0] FSM_fft_64_stage_2_0_t916;
reg [33-1:0] FSM_fft_64_stage_2_0_t917;
reg [32-1:0] FSM_fft_64_stage_2_0_t918;
reg [6-1:0] FSM_fft_64_stage_2_0_t919;
reg [32-1:0] FSM_fft_64_stage_2_0_t920;
reg [33-1:0] FSM_fft_64_stage_2_0_t921;
reg [32-1:0] FSM_fft_64_stage_2_0_t922;
reg [2048-1:0] FSM_fft_64_stage_2_0_t923;
reg [33-1:0] FSM_fft_64_stage_2_0_t924;
reg [32-1:0] FSM_fft_64_stage_2_0_t925;
reg [6-1:0] FSM_fft_64_stage_2_0_t926;
reg [2048-1:0] FSM_fft_64_stage_2_0_t927;
reg [6-1:0] FSM_fft_64_stage_2_0_t928;
reg [6-1:0] FSM_fft_64_stage_2_0_t929;
reg [32-1:0] FSM_fft_64_stage_2_0_t930;
reg [33-1:0] FSM_fft_64_stage_2_0_t931;
reg [32-1:0] FSM_fft_64_stage_2_0_t932;
reg [6-1:0] FSM_fft_64_stage_2_0_t933;
reg [32-1:0] FSM_fft_64_stage_2_0_t934;
reg [33-1:0] FSM_fft_64_stage_2_0_t935;
reg [32-1:0] FSM_fft_64_stage_2_0_t936;
reg [2048-1:0] FSM_fft_64_stage_2_0_t937;
reg [33-1:0] FSM_fft_64_stage_2_0_t938;
reg [32-1:0] FSM_fft_64_stage_2_0_t939;
reg [6-1:0] FSM_fft_64_stage_2_0_t940;
reg [2048-1:0] FSM_fft_64_stage_2_0_t941;
reg [33-1:0] FSM_fft_64_stage_2_0_t942;
reg [32-1:0] FSM_fft_64_stage_2_0_t943;
reg [6-1:0] FSM_fft_64_stage_2_0_t944;
reg [33-1:0] FSM_fft_64_stage_2_0_t945;
reg [32-1:0] FSM_fft_64_stage_2_0_t946;
reg [6-1:0] FSM_fft_64_stage_2_0_t947;
reg [32-1:0] FSM_fft_64_stage_2_0_t948;
reg [33-1:0] FSM_fft_64_stage_2_0_t949;
reg [32-1:0] FSM_fft_64_stage_2_0_t950;
reg [6-1:0] FSM_fft_64_stage_2_0_t951;
reg [32-1:0] FSM_fft_64_stage_2_0_t952;
reg [33-1:0] FSM_fft_64_stage_2_0_t953;
reg [32-1:0] FSM_fft_64_stage_2_0_t954;
reg [2048-1:0] FSM_fft_64_stage_2_0_t955;
reg [33-1:0] FSM_fft_64_stage_2_0_t956;
reg [32-1:0] FSM_fft_64_stage_2_0_t957;
reg [6-1:0] FSM_fft_64_stage_2_0_t958;
reg [2048-1:0] FSM_fft_64_stage_2_0_t959;
reg [6-1:0] FSM_fft_64_stage_2_0_t960;
reg [6-1:0] FSM_fft_64_stage_2_0_t961;
reg [32-1:0] FSM_fft_64_stage_2_0_t962;
reg [33-1:0] FSM_fft_64_stage_2_0_t963;
reg [32-1:0] FSM_fft_64_stage_2_0_t964;
reg [6-1:0] FSM_fft_64_stage_2_0_t965;
reg [32-1:0] FSM_fft_64_stage_2_0_t966;
reg [33-1:0] FSM_fft_64_stage_2_0_t967;
reg [32-1:0] FSM_fft_64_stage_2_0_t968;
reg [2048-1:0] FSM_fft_64_stage_2_0_t969;
reg [33-1:0] FSM_fft_64_stage_2_0_t970;
reg [32-1:0] FSM_fft_64_stage_2_0_t971;
reg [6-1:0] FSM_fft_64_stage_2_0_t972;
reg [2048-1:0] FSM_fft_64_stage_2_0_t973;
reg [33-1:0] FSM_fft_64_stage_2_0_t974;
reg [32-1:0] FSM_fft_64_stage_2_0_t975;
reg [6-1:0] FSM_fft_64_stage_2_0_t976;
reg [33-1:0] FSM_fft_64_stage_2_0_t977;
reg [32-1:0] FSM_fft_64_stage_2_0_t978;
reg [6-1:0] FSM_fft_64_stage_2_0_t979;
reg [32-1:0] FSM_fft_64_stage_2_0_t980;
reg [33-1:0] FSM_fft_64_stage_2_0_t981;
reg [32-1:0] FSM_fft_64_stage_2_0_t982;
reg [6-1:0] FSM_fft_64_stage_2_0_t983;
reg [32-1:0] FSM_fft_64_stage_2_0_t984;
reg [33-1:0] FSM_fft_64_stage_2_0_t985;
reg [32-1:0] FSM_fft_64_stage_2_0_t986;
reg [2048-1:0] FSM_fft_64_stage_2_0_t987;
reg [33-1:0] FSM_fft_64_stage_2_0_t988;
reg [32-1:0] FSM_fft_64_stage_2_0_t989;
reg [6-1:0] FSM_fft_64_stage_2_0_t990;
reg [2048-1:0] FSM_fft_64_stage_2_0_t991;
reg [6-1:0] FSM_fft_64_stage_2_0_t992;
reg [6-1:0] FSM_fft_64_stage_2_0_t993;
reg [32-1:0] FSM_fft_64_stage_2_0_t994;
reg [33-1:0] FSM_fft_64_stage_2_0_t995;
reg [32-1:0] FSM_fft_64_stage_2_0_t996;
reg [6-1:0] FSM_fft_64_stage_2_0_t997;
reg [32-1:0] FSM_fft_64_stage_2_0_t998;
reg [33-1:0] FSM_fft_64_stage_2_0_t999;
reg [32-1:0] FSM_fft_64_stage_2_0_t1000;
reg [2048-1:0] FSM_fft_64_stage_2_0_t1001;
reg [33-1:0] FSM_fft_64_stage_2_0_t1002;
reg [32-1:0] FSM_fft_64_stage_2_0_t1003;
reg [6-1:0] FSM_fft_64_stage_2_0_t1004;
reg [2048-1:0] FSM_fft_64_stage_2_0_t1005;
reg [33-1:0] FSM_fft_64_stage_2_0_t1006;
reg [32-1:0] FSM_fft_64_stage_2_0_t1007;
reg [6-1:0] FSM_fft_64_stage_2_0_t1008;
reg [33-1:0] FSM_fft_64_stage_2_0_t1009;
reg [32-1:0] FSM_fft_64_stage_2_0_t1010;
reg [6-1:0] FSM_fft_64_stage_2_0_t1011;
reg [32-1:0] FSM_fft_64_stage_2_0_t1012;
reg [33-1:0] FSM_fft_64_stage_2_0_t1013;
reg [32-1:0] FSM_fft_64_stage_2_0_t1014;
reg [6-1:0] FSM_fft_64_stage_2_0_t1015;
reg [32-1:0] FSM_fft_64_stage_2_0_t1016;
reg [33-1:0] FSM_fft_64_stage_2_0_t1017;
reg [32-1:0] FSM_fft_64_stage_2_0_t1018;
reg [2048-1:0] FSM_fft_64_stage_2_0_t1019;
reg [33-1:0] FSM_fft_64_stage_2_0_t1020;
reg [32-1:0] FSM_fft_64_stage_2_0_t1021;
reg [6-1:0] FSM_fft_64_stage_2_0_t1022;
reg [2048-1:0] FSM_fft_64_stage_2_0_t1023;
reg [6-1:0] FSM_fft_64_stage_2_0_t1024;
reg [6-1:0] FSM_fft_64_stage_2_0_t1025;
reg [32-1:0] FSM_fft_64_stage_2_0_t1026;
reg [33-1:0] FSM_fft_64_stage_2_0_t1027;
reg [32-1:0] FSM_fft_64_stage_2_0_t1028;
reg [6-1:0] FSM_fft_64_stage_2_0_t1029;
reg [32-1:0] FSM_fft_64_stage_2_0_t1030;
reg [33-1:0] FSM_fft_64_stage_2_0_t1031;
reg [32-1:0] FSM_fft_64_stage_2_0_t1032;
reg [2048-1:0] FSM_fft_64_stage_2_0_t1033;
reg [33-1:0] FSM_fft_64_stage_2_0_t1034;
reg [32-1:0] FSM_fft_64_stage_2_0_t1035;
reg [6-1:0] FSM_fft_64_stage_2_0_t1036;
reg [2048-1:0] FSM_fft_64_stage_2_0_t1037;
reg [33-1:0] FSM_fft_64_stage_2_0_t1038;
reg [32-1:0] FSM_fft_64_stage_2_0_t1039;
reg [6-1:0] FSM_fft_64_stage_2_0_t1040;
reg [33-1:0] FSM_fft_64_stage_2_0_t1041;
reg [32-1:0] FSM_fft_64_stage_2_0_t1042;
reg [6-1:0] FSM_fft_64_stage_2_0_t1043;
reg [32-1:0] FSM_fft_64_stage_2_0_t1044;
reg [33-1:0] FSM_fft_64_stage_2_0_t1045;
reg [32-1:0] FSM_fft_64_stage_2_0_t1046;
reg [6-1:0] FSM_fft_64_stage_2_0_t1047;
reg [32-1:0] FSM_fft_64_stage_2_0_t1048;
reg [33-1:0] FSM_fft_64_stage_2_0_t1049;
reg [32-1:0] FSM_fft_64_stage_2_0_t1050;
reg [2048-1:0] FSM_fft_64_stage_2_0_t1051;
reg [33-1:0] FSM_fft_64_stage_2_0_t1052;
reg [32-1:0] FSM_fft_64_stage_2_0_t1053;
reg [6-1:0] FSM_fft_64_stage_2_0_t1054;
reg [2048-1:0] FSM_fft_64_stage_2_0_t1055;

assign FSM_fft_64_stage_2_0_out_valid = 1'b1;
/*
    Wiring by fft_64_stage_2
*/
assign i_ready = FSM_fft_64_stage_2_0_in_ready;
assign o_data_out_real = FSM_fft_64_stage_2_0_t543;
assign o_data_out_imag = FSM_fft_64_stage_2_0_t1055;
assign o_valid = FSM_fft_64_stage_2_0_out_valid;
/* End wiring by fft_64_stage_2 */

initial begin
    FSM_fft_64_stage_2_0_t0 = 32'b0 * 32'b00000000000000000000000000000100;
    FSM_fft_64_stage_2_0_t1 = FSM_fft_64_stage_2_0_t0[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t2 = FSM_fft_64_stage_2_0_t1[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t3 = FSM_fft_64_stage_2_0_t1[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t4 = i_data_in_real[FSM_fft_64_stage_2_0_t3 * 32 +: 32];
    FSM_fft_64_stage_2_0_t5 = FSM_fft_64_stage_2_0_t1 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t6 = FSM_fft_64_stage_2_0_t5[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t7 = FSM_fft_64_stage_2_0_t6[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t8 = i_data_in_real[FSM_fft_64_stage_2_0_t7 * 32 +: 32];
    FSM_fft_64_stage_2_0_t9 = FSM_fft_64_stage_2_0_t4 + FSM_fft_64_stage_2_0_t8;
    FSM_fft_64_stage_2_0_t10 = FSM_fft_64_stage_2_0_t9[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t11 = i_data_in_real;
    FSM_fft_64_stage_2_0_t11[FSM_fft_64_stage_2_0_t2 * 32 +: 32] = FSM_fft_64_stage_2_0_t10;
    FSM_fft_64_stage_2_0_t12 = FSM_fft_64_stage_2_0_t1 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t13 = FSM_fft_64_stage_2_0_t12[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t14 = FSM_fft_64_stage_2_0_t13[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t15 = FSM_fft_64_stage_2_0_t11;
    FSM_fft_64_stage_2_0_t15[FSM_fft_64_stage_2_0_t14 * 32 +: 32] = FSM_fft_64_stage_2_0_t4 - FSM_fft_64_stage_2_0_t8;
    FSM_fft_64_stage_2_0_t16 = FSM_fft_64_stage_2_0_t1 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t17 = FSM_fft_64_stage_2_0_t16[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t18 = FSM_fft_64_stage_2_0_t17[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t19 = FSM_fft_64_stage_2_0_t1 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t20 = FSM_fft_64_stage_2_0_t19[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t21 = FSM_fft_64_stage_2_0_t20[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t22 = i_data_in_real[FSM_fft_64_stage_2_0_t21 * 32 +: 32];
    FSM_fft_64_stage_2_0_t23 = FSM_fft_64_stage_2_0_t1 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t24 = FSM_fft_64_stage_2_0_t23[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t25 = FSM_fft_64_stage_2_0_t24[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t26 = i_data_in_real[FSM_fft_64_stage_2_0_t25 * 32 +: 32];
    FSM_fft_64_stage_2_0_t27 = FSM_fft_64_stage_2_0_t22 + FSM_fft_64_stage_2_0_t26;
    FSM_fft_64_stage_2_0_t28 = FSM_fft_64_stage_2_0_t27[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t29 = FSM_fft_64_stage_2_0_t15;
    FSM_fft_64_stage_2_0_t29[FSM_fft_64_stage_2_0_t18 * 32 +: 32] = FSM_fft_64_stage_2_0_t28;
    FSM_fft_64_stage_2_0_t30 = FSM_fft_64_stage_2_0_t1 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t31 = FSM_fft_64_stage_2_0_t30[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t32 = FSM_fft_64_stage_2_0_t31[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t33 = FSM_fft_64_stage_2_0_t29;
    FSM_fft_64_stage_2_0_t33[FSM_fft_64_stage_2_0_t32 * 32 +: 32] = FSM_fft_64_stage_2_0_t22 - FSM_fft_64_stage_2_0_t26;
    FSM_fft_64_stage_2_0_t34 = 32'b00000000000000000000000000000001 * 32'b00000000000000000000000000000100;
    FSM_fft_64_stage_2_0_t35 = FSM_fft_64_stage_2_0_t34[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t36 = FSM_fft_64_stage_2_0_t35[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t37 = FSM_fft_64_stage_2_0_t35[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t38 = FSM_fft_64_stage_2_0_t33[FSM_fft_64_stage_2_0_t37 * 32 +: 32];
    FSM_fft_64_stage_2_0_t39 = FSM_fft_64_stage_2_0_t35 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t40 = FSM_fft_64_stage_2_0_t39[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t41 = FSM_fft_64_stage_2_0_t40[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t42 = FSM_fft_64_stage_2_0_t33[FSM_fft_64_stage_2_0_t41 * 32 +: 32];
    FSM_fft_64_stage_2_0_t43 = FSM_fft_64_stage_2_0_t38 + FSM_fft_64_stage_2_0_t42;
    FSM_fft_64_stage_2_0_t44 = FSM_fft_64_stage_2_0_t43[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t45 = FSM_fft_64_stage_2_0_t33;
    FSM_fft_64_stage_2_0_t45[FSM_fft_64_stage_2_0_t36 * 32 +: 32] = FSM_fft_64_stage_2_0_t44;
    FSM_fft_64_stage_2_0_t46 = FSM_fft_64_stage_2_0_t35 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t47 = FSM_fft_64_stage_2_0_t46[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t48 = FSM_fft_64_stage_2_0_t47[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t49 = FSM_fft_64_stage_2_0_t45;
    FSM_fft_64_stage_2_0_t49[FSM_fft_64_stage_2_0_t48 * 32 +: 32] = FSM_fft_64_stage_2_0_t38 - FSM_fft_64_stage_2_0_t42;
    FSM_fft_64_stage_2_0_t50 = FSM_fft_64_stage_2_0_t35 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t51 = FSM_fft_64_stage_2_0_t50[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t52 = FSM_fft_64_stage_2_0_t51[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t53 = FSM_fft_64_stage_2_0_t35 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t54 = FSM_fft_64_stage_2_0_t53[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t55 = FSM_fft_64_stage_2_0_t54[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t56 = FSM_fft_64_stage_2_0_t33[FSM_fft_64_stage_2_0_t55 * 32 +: 32];
    FSM_fft_64_stage_2_0_t57 = FSM_fft_64_stage_2_0_t35 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t58 = FSM_fft_64_stage_2_0_t57[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t59 = FSM_fft_64_stage_2_0_t58[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t60 = FSM_fft_64_stage_2_0_t33[FSM_fft_64_stage_2_0_t59 * 32 +: 32];
    FSM_fft_64_stage_2_0_t61 = FSM_fft_64_stage_2_0_t56 + FSM_fft_64_stage_2_0_t60;
    FSM_fft_64_stage_2_0_t62 = FSM_fft_64_stage_2_0_t61[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t63 = FSM_fft_64_stage_2_0_t49;
    FSM_fft_64_stage_2_0_t63[FSM_fft_64_stage_2_0_t52 * 32 +: 32] = FSM_fft_64_stage_2_0_t62;
    FSM_fft_64_stage_2_0_t64 = FSM_fft_64_stage_2_0_t35 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t65 = FSM_fft_64_stage_2_0_t64[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t66 = FSM_fft_64_stage_2_0_t65[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t67 = FSM_fft_64_stage_2_0_t63;
    FSM_fft_64_stage_2_0_t67[FSM_fft_64_stage_2_0_t66 * 32 +: 32] = FSM_fft_64_stage_2_0_t56 - FSM_fft_64_stage_2_0_t60;
    FSM_fft_64_stage_2_0_t68 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000100;
    FSM_fft_64_stage_2_0_t69 = FSM_fft_64_stage_2_0_t68[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t70 = FSM_fft_64_stage_2_0_t69[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t71 = FSM_fft_64_stage_2_0_t69[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t72 = FSM_fft_64_stage_2_0_t67[FSM_fft_64_stage_2_0_t71 * 32 +: 32];
    FSM_fft_64_stage_2_0_t73 = FSM_fft_64_stage_2_0_t69 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t74 = FSM_fft_64_stage_2_0_t73[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t75 = FSM_fft_64_stage_2_0_t74[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t76 = FSM_fft_64_stage_2_0_t67[FSM_fft_64_stage_2_0_t75 * 32 +: 32];
    FSM_fft_64_stage_2_0_t77 = FSM_fft_64_stage_2_0_t72 + FSM_fft_64_stage_2_0_t76;
    FSM_fft_64_stage_2_0_t78 = FSM_fft_64_stage_2_0_t77[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t79 = FSM_fft_64_stage_2_0_t67;
    FSM_fft_64_stage_2_0_t79[FSM_fft_64_stage_2_0_t70 * 32 +: 32] = FSM_fft_64_stage_2_0_t78;
    FSM_fft_64_stage_2_0_t80 = FSM_fft_64_stage_2_0_t69 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t81 = FSM_fft_64_stage_2_0_t80[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t82 = FSM_fft_64_stage_2_0_t81[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t83 = FSM_fft_64_stage_2_0_t79;
    FSM_fft_64_stage_2_0_t83[FSM_fft_64_stage_2_0_t82 * 32 +: 32] = FSM_fft_64_stage_2_0_t72 - FSM_fft_64_stage_2_0_t76;
    FSM_fft_64_stage_2_0_t84 = FSM_fft_64_stage_2_0_t69 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t85 = FSM_fft_64_stage_2_0_t84[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t86 = FSM_fft_64_stage_2_0_t85[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t87 = FSM_fft_64_stage_2_0_t69 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t88 = FSM_fft_64_stage_2_0_t87[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t89 = FSM_fft_64_stage_2_0_t88[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t90 = FSM_fft_64_stage_2_0_t67[FSM_fft_64_stage_2_0_t89 * 32 +: 32];
    FSM_fft_64_stage_2_0_t91 = FSM_fft_64_stage_2_0_t69 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t92 = FSM_fft_64_stage_2_0_t91[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t93 = FSM_fft_64_stage_2_0_t92[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t94 = FSM_fft_64_stage_2_0_t67[FSM_fft_64_stage_2_0_t93 * 32 +: 32];
    FSM_fft_64_stage_2_0_t95 = FSM_fft_64_stage_2_0_t90 + FSM_fft_64_stage_2_0_t94;
    FSM_fft_64_stage_2_0_t96 = FSM_fft_64_stage_2_0_t95[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t97 = FSM_fft_64_stage_2_0_t83;
    FSM_fft_64_stage_2_0_t97[FSM_fft_64_stage_2_0_t86 * 32 +: 32] = FSM_fft_64_stage_2_0_t96;
    FSM_fft_64_stage_2_0_t98 = FSM_fft_64_stage_2_0_t69 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t99 = FSM_fft_64_stage_2_0_t98[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t100 = FSM_fft_64_stage_2_0_t99[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t101 = FSM_fft_64_stage_2_0_t97;
    FSM_fft_64_stage_2_0_t101[FSM_fft_64_stage_2_0_t100 * 32 +: 32] = FSM_fft_64_stage_2_0_t90 - FSM_fft_64_stage_2_0_t94;
    FSM_fft_64_stage_2_0_t102 = 32'b00000000000000000000000000000011 * 32'b00000000000000000000000000000100;
    FSM_fft_64_stage_2_0_t103 = FSM_fft_64_stage_2_0_t102[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t104 = FSM_fft_64_stage_2_0_t103[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t105 = FSM_fft_64_stage_2_0_t103[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t106 = FSM_fft_64_stage_2_0_t101[FSM_fft_64_stage_2_0_t105 * 32 +: 32];
    FSM_fft_64_stage_2_0_t107 = FSM_fft_64_stage_2_0_t103 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t108 = FSM_fft_64_stage_2_0_t107[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t109 = FSM_fft_64_stage_2_0_t108[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t110 = FSM_fft_64_stage_2_0_t101[FSM_fft_64_stage_2_0_t109 * 32 +: 32];
    FSM_fft_64_stage_2_0_t111 = FSM_fft_64_stage_2_0_t106 + FSM_fft_64_stage_2_0_t110;
    FSM_fft_64_stage_2_0_t112 = FSM_fft_64_stage_2_0_t111[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t113 = FSM_fft_64_stage_2_0_t101;
    FSM_fft_64_stage_2_0_t113[FSM_fft_64_stage_2_0_t104 * 32 +: 32] = FSM_fft_64_stage_2_0_t112;
    FSM_fft_64_stage_2_0_t114 = FSM_fft_64_stage_2_0_t103 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t115 = FSM_fft_64_stage_2_0_t114[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t116 = FSM_fft_64_stage_2_0_t115[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t117 = FSM_fft_64_stage_2_0_t113;
    FSM_fft_64_stage_2_0_t117[FSM_fft_64_stage_2_0_t116 * 32 +: 32] = FSM_fft_64_stage_2_0_t106 - FSM_fft_64_stage_2_0_t110;
    FSM_fft_64_stage_2_0_t118 = FSM_fft_64_stage_2_0_t103 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t119 = FSM_fft_64_stage_2_0_t118[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t120 = FSM_fft_64_stage_2_0_t119[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t121 = FSM_fft_64_stage_2_0_t103 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t122 = FSM_fft_64_stage_2_0_t121[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t123 = FSM_fft_64_stage_2_0_t122[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t124 = FSM_fft_64_stage_2_0_t101[FSM_fft_64_stage_2_0_t123 * 32 +: 32];
    FSM_fft_64_stage_2_0_t125 = FSM_fft_64_stage_2_0_t103 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t126 = FSM_fft_64_stage_2_0_t125[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t127 = FSM_fft_64_stage_2_0_t126[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t128 = FSM_fft_64_stage_2_0_t101[FSM_fft_64_stage_2_0_t127 * 32 +: 32];
    FSM_fft_64_stage_2_0_t129 = FSM_fft_64_stage_2_0_t124 + FSM_fft_64_stage_2_0_t128;
    FSM_fft_64_stage_2_0_t130 = FSM_fft_64_stage_2_0_t129[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t131 = FSM_fft_64_stage_2_0_t117;
    FSM_fft_64_stage_2_0_t131[FSM_fft_64_stage_2_0_t120 * 32 +: 32] = FSM_fft_64_stage_2_0_t130;
    FSM_fft_64_stage_2_0_t132 = FSM_fft_64_stage_2_0_t103 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t133 = FSM_fft_64_stage_2_0_t132[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t134 = FSM_fft_64_stage_2_0_t133[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t135 = FSM_fft_64_stage_2_0_t131;
    FSM_fft_64_stage_2_0_t135[FSM_fft_64_stage_2_0_t134 * 32 +: 32] = FSM_fft_64_stage_2_0_t124 - FSM_fft_64_stage_2_0_t128;
    FSM_fft_64_stage_2_0_t136 = 32'b00000000000000000000000000000100 * 32'b00000000000000000000000000000100;
    FSM_fft_64_stage_2_0_t137 = FSM_fft_64_stage_2_0_t136[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t138 = FSM_fft_64_stage_2_0_t137[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t139 = FSM_fft_64_stage_2_0_t137[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t140 = FSM_fft_64_stage_2_0_t135[FSM_fft_64_stage_2_0_t139 * 32 +: 32];
    FSM_fft_64_stage_2_0_t141 = FSM_fft_64_stage_2_0_t137 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t142 = FSM_fft_64_stage_2_0_t141[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t143 = FSM_fft_64_stage_2_0_t142[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t144 = FSM_fft_64_stage_2_0_t135[FSM_fft_64_stage_2_0_t143 * 32 +: 32];
    FSM_fft_64_stage_2_0_t145 = FSM_fft_64_stage_2_0_t140 + FSM_fft_64_stage_2_0_t144;
    FSM_fft_64_stage_2_0_t146 = FSM_fft_64_stage_2_0_t145[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t147 = FSM_fft_64_stage_2_0_t135;
    FSM_fft_64_stage_2_0_t147[FSM_fft_64_stage_2_0_t138 * 32 +: 32] = FSM_fft_64_stage_2_0_t146;
    FSM_fft_64_stage_2_0_t148 = FSM_fft_64_stage_2_0_t137 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t149 = FSM_fft_64_stage_2_0_t148[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t150 = FSM_fft_64_stage_2_0_t149[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t151 = FSM_fft_64_stage_2_0_t147;
    FSM_fft_64_stage_2_0_t151[FSM_fft_64_stage_2_0_t150 * 32 +: 32] = FSM_fft_64_stage_2_0_t140 - FSM_fft_64_stage_2_0_t144;
    FSM_fft_64_stage_2_0_t152 = FSM_fft_64_stage_2_0_t137 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t153 = FSM_fft_64_stage_2_0_t152[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t154 = FSM_fft_64_stage_2_0_t153[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t155 = FSM_fft_64_stage_2_0_t137 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t156 = FSM_fft_64_stage_2_0_t155[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t157 = FSM_fft_64_stage_2_0_t156[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t158 = FSM_fft_64_stage_2_0_t135[FSM_fft_64_stage_2_0_t157 * 32 +: 32];
    FSM_fft_64_stage_2_0_t159 = FSM_fft_64_stage_2_0_t137 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t160 = FSM_fft_64_stage_2_0_t159[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t161 = FSM_fft_64_stage_2_0_t160[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t162 = FSM_fft_64_stage_2_0_t135[FSM_fft_64_stage_2_0_t161 * 32 +: 32];
    FSM_fft_64_stage_2_0_t163 = FSM_fft_64_stage_2_0_t158 + FSM_fft_64_stage_2_0_t162;
    FSM_fft_64_stage_2_0_t164 = FSM_fft_64_stage_2_0_t163[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t165 = FSM_fft_64_stage_2_0_t151;
    FSM_fft_64_stage_2_0_t165[FSM_fft_64_stage_2_0_t154 * 32 +: 32] = FSM_fft_64_stage_2_0_t164;
    FSM_fft_64_stage_2_0_t166 = FSM_fft_64_stage_2_0_t137 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t167 = FSM_fft_64_stage_2_0_t166[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t168 = FSM_fft_64_stage_2_0_t167[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t169 = FSM_fft_64_stage_2_0_t165;
    FSM_fft_64_stage_2_0_t169[FSM_fft_64_stage_2_0_t168 * 32 +: 32] = FSM_fft_64_stage_2_0_t158 - FSM_fft_64_stage_2_0_t162;
    FSM_fft_64_stage_2_0_t170 = 32'b00000000000000000000000000000101 * 32'b00000000000000000000000000000100;
    FSM_fft_64_stage_2_0_t171 = FSM_fft_64_stage_2_0_t170[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t172 = FSM_fft_64_stage_2_0_t171[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t173 = FSM_fft_64_stage_2_0_t171[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t174 = FSM_fft_64_stage_2_0_t169[FSM_fft_64_stage_2_0_t173 * 32 +: 32];
    FSM_fft_64_stage_2_0_t175 = FSM_fft_64_stage_2_0_t171 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t176 = FSM_fft_64_stage_2_0_t175[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t177 = FSM_fft_64_stage_2_0_t176[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t178 = FSM_fft_64_stage_2_0_t169[FSM_fft_64_stage_2_0_t177 * 32 +: 32];
    FSM_fft_64_stage_2_0_t179 = FSM_fft_64_stage_2_0_t174 + FSM_fft_64_stage_2_0_t178;
    FSM_fft_64_stage_2_0_t180 = FSM_fft_64_stage_2_0_t179[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t181 = FSM_fft_64_stage_2_0_t169;
    FSM_fft_64_stage_2_0_t181[FSM_fft_64_stage_2_0_t172 * 32 +: 32] = FSM_fft_64_stage_2_0_t180;
    FSM_fft_64_stage_2_0_t182 = FSM_fft_64_stage_2_0_t171 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t183 = FSM_fft_64_stage_2_0_t182[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t184 = FSM_fft_64_stage_2_0_t183[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t185 = FSM_fft_64_stage_2_0_t181;
    FSM_fft_64_stage_2_0_t185[FSM_fft_64_stage_2_0_t184 * 32 +: 32] = FSM_fft_64_stage_2_0_t174 - FSM_fft_64_stage_2_0_t178;
    FSM_fft_64_stage_2_0_t186 = FSM_fft_64_stage_2_0_t171 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t187 = FSM_fft_64_stage_2_0_t186[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t188 = FSM_fft_64_stage_2_0_t187[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t189 = FSM_fft_64_stage_2_0_t171 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t190 = FSM_fft_64_stage_2_0_t189[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t191 = FSM_fft_64_stage_2_0_t190[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t192 = FSM_fft_64_stage_2_0_t169[FSM_fft_64_stage_2_0_t191 * 32 +: 32];
    FSM_fft_64_stage_2_0_t193 = FSM_fft_64_stage_2_0_t171 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t194 = FSM_fft_64_stage_2_0_t193[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t195 = FSM_fft_64_stage_2_0_t194[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t196 = FSM_fft_64_stage_2_0_t169[FSM_fft_64_stage_2_0_t195 * 32 +: 32];
    FSM_fft_64_stage_2_0_t197 = FSM_fft_64_stage_2_0_t192 + FSM_fft_64_stage_2_0_t196;
    FSM_fft_64_stage_2_0_t198 = FSM_fft_64_stage_2_0_t197[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t199 = FSM_fft_64_stage_2_0_t185;
    FSM_fft_64_stage_2_0_t199[FSM_fft_64_stage_2_0_t188 * 32 +: 32] = FSM_fft_64_stage_2_0_t198;
    FSM_fft_64_stage_2_0_t200 = FSM_fft_64_stage_2_0_t171 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t201 = FSM_fft_64_stage_2_0_t200[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t202 = FSM_fft_64_stage_2_0_t201[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t203 = FSM_fft_64_stage_2_0_t199;
    FSM_fft_64_stage_2_0_t203[FSM_fft_64_stage_2_0_t202 * 32 +: 32] = FSM_fft_64_stage_2_0_t192 - FSM_fft_64_stage_2_0_t196;
    FSM_fft_64_stage_2_0_t204 = 32'b00000000000000000000000000000110 * 32'b00000000000000000000000000000100;
    FSM_fft_64_stage_2_0_t205 = FSM_fft_64_stage_2_0_t204[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t206 = FSM_fft_64_stage_2_0_t205[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t207 = FSM_fft_64_stage_2_0_t205[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t208 = FSM_fft_64_stage_2_0_t203[FSM_fft_64_stage_2_0_t207 * 32 +: 32];
    FSM_fft_64_stage_2_0_t209 = FSM_fft_64_stage_2_0_t205 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t210 = FSM_fft_64_stage_2_0_t209[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t211 = FSM_fft_64_stage_2_0_t210[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t212 = FSM_fft_64_stage_2_0_t203[FSM_fft_64_stage_2_0_t211 * 32 +: 32];
    FSM_fft_64_stage_2_0_t213 = FSM_fft_64_stage_2_0_t208 + FSM_fft_64_stage_2_0_t212;
    FSM_fft_64_stage_2_0_t214 = FSM_fft_64_stage_2_0_t213[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t215 = FSM_fft_64_stage_2_0_t203;
    FSM_fft_64_stage_2_0_t215[FSM_fft_64_stage_2_0_t206 * 32 +: 32] = FSM_fft_64_stage_2_0_t214;
    FSM_fft_64_stage_2_0_t216 = FSM_fft_64_stage_2_0_t205 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t217 = FSM_fft_64_stage_2_0_t216[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t218 = FSM_fft_64_stage_2_0_t217[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t219 = FSM_fft_64_stage_2_0_t215;
    FSM_fft_64_stage_2_0_t219[FSM_fft_64_stage_2_0_t218 * 32 +: 32] = FSM_fft_64_stage_2_0_t208 - FSM_fft_64_stage_2_0_t212;
    FSM_fft_64_stage_2_0_t220 = FSM_fft_64_stage_2_0_t205 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t221 = FSM_fft_64_stage_2_0_t220[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t222 = FSM_fft_64_stage_2_0_t221[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t223 = FSM_fft_64_stage_2_0_t205 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t224 = FSM_fft_64_stage_2_0_t223[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t225 = FSM_fft_64_stage_2_0_t224[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t226 = FSM_fft_64_stage_2_0_t203[FSM_fft_64_stage_2_0_t225 * 32 +: 32];
    FSM_fft_64_stage_2_0_t227 = FSM_fft_64_stage_2_0_t205 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t228 = FSM_fft_64_stage_2_0_t227[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t229 = FSM_fft_64_stage_2_0_t228[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t230 = FSM_fft_64_stage_2_0_t203[FSM_fft_64_stage_2_0_t229 * 32 +: 32];
    FSM_fft_64_stage_2_0_t231 = FSM_fft_64_stage_2_0_t226 + FSM_fft_64_stage_2_0_t230;
    FSM_fft_64_stage_2_0_t232 = FSM_fft_64_stage_2_0_t231[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t233 = FSM_fft_64_stage_2_0_t219;
    FSM_fft_64_stage_2_0_t233[FSM_fft_64_stage_2_0_t222 * 32 +: 32] = FSM_fft_64_stage_2_0_t232;
    FSM_fft_64_stage_2_0_t234 = FSM_fft_64_stage_2_0_t205 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t235 = FSM_fft_64_stage_2_0_t234[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t236 = FSM_fft_64_stage_2_0_t235[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t237 = FSM_fft_64_stage_2_0_t233;
    FSM_fft_64_stage_2_0_t237[FSM_fft_64_stage_2_0_t236 * 32 +: 32] = FSM_fft_64_stage_2_0_t226 - FSM_fft_64_stage_2_0_t230;
    FSM_fft_64_stage_2_0_t238 = 32'b00000000000000000000000000000111 * 32'b00000000000000000000000000000100;
    FSM_fft_64_stage_2_0_t239 = FSM_fft_64_stage_2_0_t238[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t240 = FSM_fft_64_stage_2_0_t239[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t241 = FSM_fft_64_stage_2_0_t239[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t242 = FSM_fft_64_stage_2_0_t237[FSM_fft_64_stage_2_0_t241 * 32 +: 32];
    FSM_fft_64_stage_2_0_t243 = FSM_fft_64_stage_2_0_t239 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t244 = FSM_fft_64_stage_2_0_t243[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t245 = FSM_fft_64_stage_2_0_t244[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t246 = FSM_fft_64_stage_2_0_t237[FSM_fft_64_stage_2_0_t245 * 32 +: 32];
    FSM_fft_64_stage_2_0_t247 = FSM_fft_64_stage_2_0_t242 + FSM_fft_64_stage_2_0_t246;
    FSM_fft_64_stage_2_0_t248 = FSM_fft_64_stage_2_0_t247[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t249 = FSM_fft_64_stage_2_0_t237;
    FSM_fft_64_stage_2_0_t249[FSM_fft_64_stage_2_0_t240 * 32 +: 32] = FSM_fft_64_stage_2_0_t248;
    FSM_fft_64_stage_2_0_t250 = FSM_fft_64_stage_2_0_t239 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t251 = FSM_fft_64_stage_2_0_t250[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t252 = FSM_fft_64_stage_2_0_t251[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t253 = FSM_fft_64_stage_2_0_t249;
    FSM_fft_64_stage_2_0_t253[FSM_fft_64_stage_2_0_t252 * 32 +: 32] = FSM_fft_64_stage_2_0_t242 - FSM_fft_64_stage_2_0_t246;
    FSM_fft_64_stage_2_0_t254 = FSM_fft_64_stage_2_0_t239 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t255 = FSM_fft_64_stage_2_0_t254[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t256 = FSM_fft_64_stage_2_0_t255[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t257 = FSM_fft_64_stage_2_0_t239 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t258 = FSM_fft_64_stage_2_0_t257[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t259 = FSM_fft_64_stage_2_0_t258[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t260 = FSM_fft_64_stage_2_0_t237[FSM_fft_64_stage_2_0_t259 * 32 +: 32];
    FSM_fft_64_stage_2_0_t261 = FSM_fft_64_stage_2_0_t239 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t262 = FSM_fft_64_stage_2_0_t261[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t263 = FSM_fft_64_stage_2_0_t262[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t264 = FSM_fft_64_stage_2_0_t237[FSM_fft_64_stage_2_0_t263 * 32 +: 32];
    FSM_fft_64_stage_2_0_t265 = FSM_fft_64_stage_2_0_t260 + FSM_fft_64_stage_2_0_t264;
    FSM_fft_64_stage_2_0_t266 = FSM_fft_64_stage_2_0_t265[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t267 = FSM_fft_64_stage_2_0_t253;
    FSM_fft_64_stage_2_0_t267[FSM_fft_64_stage_2_0_t256 * 32 +: 32] = FSM_fft_64_stage_2_0_t266;
    FSM_fft_64_stage_2_0_t268 = FSM_fft_64_stage_2_0_t239 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t269 = FSM_fft_64_stage_2_0_t268[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t270 = FSM_fft_64_stage_2_0_t269[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t271 = FSM_fft_64_stage_2_0_t267;
    FSM_fft_64_stage_2_0_t271[FSM_fft_64_stage_2_0_t270 * 32 +: 32] = FSM_fft_64_stage_2_0_t260 - FSM_fft_64_stage_2_0_t264;
    FSM_fft_64_stage_2_0_t272 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_fft_64_stage_2_0_t273 = FSM_fft_64_stage_2_0_t272[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t274 = FSM_fft_64_stage_2_0_t273[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t275 = FSM_fft_64_stage_2_0_t273[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t276 = FSM_fft_64_stage_2_0_t271[FSM_fft_64_stage_2_0_t275 * 32 +: 32];
    FSM_fft_64_stage_2_0_t277 = FSM_fft_64_stage_2_0_t273 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t278 = FSM_fft_64_stage_2_0_t277[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t279 = FSM_fft_64_stage_2_0_t278[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t280 = FSM_fft_64_stage_2_0_t271[FSM_fft_64_stage_2_0_t279 * 32 +: 32];
    FSM_fft_64_stage_2_0_t281 = FSM_fft_64_stage_2_0_t276 + FSM_fft_64_stage_2_0_t280;
    FSM_fft_64_stage_2_0_t282 = FSM_fft_64_stage_2_0_t281[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t283 = FSM_fft_64_stage_2_0_t271;
    FSM_fft_64_stage_2_0_t283[FSM_fft_64_stage_2_0_t274 * 32 +: 32] = FSM_fft_64_stage_2_0_t282;
    FSM_fft_64_stage_2_0_t284 = FSM_fft_64_stage_2_0_t273 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t285 = FSM_fft_64_stage_2_0_t284[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t286 = FSM_fft_64_stage_2_0_t285[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t287 = FSM_fft_64_stage_2_0_t283;
    FSM_fft_64_stage_2_0_t287[FSM_fft_64_stage_2_0_t286 * 32 +: 32] = FSM_fft_64_stage_2_0_t276 - FSM_fft_64_stage_2_0_t280;
    FSM_fft_64_stage_2_0_t288 = FSM_fft_64_stage_2_0_t273 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t289 = FSM_fft_64_stage_2_0_t288[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t290 = FSM_fft_64_stage_2_0_t289[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t291 = FSM_fft_64_stage_2_0_t273 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t292 = FSM_fft_64_stage_2_0_t291[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t293 = FSM_fft_64_stage_2_0_t292[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t294 = FSM_fft_64_stage_2_0_t271[FSM_fft_64_stage_2_0_t293 * 32 +: 32];
    FSM_fft_64_stage_2_0_t295 = FSM_fft_64_stage_2_0_t273 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t296 = FSM_fft_64_stage_2_0_t295[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t297 = FSM_fft_64_stage_2_0_t296[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t298 = FSM_fft_64_stage_2_0_t271[FSM_fft_64_stage_2_0_t297 * 32 +: 32];
    FSM_fft_64_stage_2_0_t299 = FSM_fft_64_stage_2_0_t294 + FSM_fft_64_stage_2_0_t298;
    FSM_fft_64_stage_2_0_t300 = FSM_fft_64_stage_2_0_t299[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t301 = FSM_fft_64_stage_2_0_t287;
    FSM_fft_64_stage_2_0_t301[FSM_fft_64_stage_2_0_t290 * 32 +: 32] = FSM_fft_64_stage_2_0_t300;
    FSM_fft_64_stage_2_0_t302 = FSM_fft_64_stage_2_0_t273 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t303 = FSM_fft_64_stage_2_0_t302[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t304 = FSM_fft_64_stage_2_0_t303[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t305 = FSM_fft_64_stage_2_0_t301;
    FSM_fft_64_stage_2_0_t305[FSM_fft_64_stage_2_0_t304 * 32 +: 32] = FSM_fft_64_stage_2_0_t294 - FSM_fft_64_stage_2_0_t298;
    FSM_fft_64_stage_2_0_t306 = 32'b00000000000000000000000000001001 * 32'b00000000000000000000000000000100;
    FSM_fft_64_stage_2_0_t307 = FSM_fft_64_stage_2_0_t306[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t308 = FSM_fft_64_stage_2_0_t307[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t309 = FSM_fft_64_stage_2_0_t307[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t310 = FSM_fft_64_stage_2_0_t305[FSM_fft_64_stage_2_0_t309 * 32 +: 32];
    FSM_fft_64_stage_2_0_t311 = FSM_fft_64_stage_2_0_t307 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t312 = FSM_fft_64_stage_2_0_t311[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t313 = FSM_fft_64_stage_2_0_t312[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t314 = FSM_fft_64_stage_2_0_t305[FSM_fft_64_stage_2_0_t313 * 32 +: 32];
    FSM_fft_64_stage_2_0_t315 = FSM_fft_64_stage_2_0_t310 + FSM_fft_64_stage_2_0_t314;
    FSM_fft_64_stage_2_0_t316 = FSM_fft_64_stage_2_0_t315[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t317 = FSM_fft_64_stage_2_0_t305;
    FSM_fft_64_stage_2_0_t317[FSM_fft_64_stage_2_0_t308 * 32 +: 32] = FSM_fft_64_stage_2_0_t316;
    FSM_fft_64_stage_2_0_t318 = FSM_fft_64_stage_2_0_t307 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t319 = FSM_fft_64_stage_2_0_t318[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t320 = FSM_fft_64_stage_2_0_t319[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t321 = FSM_fft_64_stage_2_0_t317;
    FSM_fft_64_stage_2_0_t321[FSM_fft_64_stage_2_0_t320 * 32 +: 32] = FSM_fft_64_stage_2_0_t310 - FSM_fft_64_stage_2_0_t314;
    FSM_fft_64_stage_2_0_t322 = FSM_fft_64_stage_2_0_t307 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t323 = FSM_fft_64_stage_2_0_t322[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t324 = FSM_fft_64_stage_2_0_t323[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t325 = FSM_fft_64_stage_2_0_t307 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t326 = FSM_fft_64_stage_2_0_t325[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t327 = FSM_fft_64_stage_2_0_t326[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t328 = FSM_fft_64_stage_2_0_t305[FSM_fft_64_stage_2_0_t327 * 32 +: 32];
    FSM_fft_64_stage_2_0_t329 = FSM_fft_64_stage_2_0_t307 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t330 = FSM_fft_64_stage_2_0_t329[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t331 = FSM_fft_64_stage_2_0_t330[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t332 = FSM_fft_64_stage_2_0_t305[FSM_fft_64_stage_2_0_t331 * 32 +: 32];
    FSM_fft_64_stage_2_0_t333 = FSM_fft_64_stage_2_0_t328 + FSM_fft_64_stage_2_0_t332;
    FSM_fft_64_stage_2_0_t334 = FSM_fft_64_stage_2_0_t333[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t335 = FSM_fft_64_stage_2_0_t321;
    FSM_fft_64_stage_2_0_t335[FSM_fft_64_stage_2_0_t324 * 32 +: 32] = FSM_fft_64_stage_2_0_t334;
    FSM_fft_64_stage_2_0_t336 = FSM_fft_64_stage_2_0_t307 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t337 = FSM_fft_64_stage_2_0_t336[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t338 = FSM_fft_64_stage_2_0_t337[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t339 = FSM_fft_64_stage_2_0_t335;
    FSM_fft_64_stage_2_0_t339[FSM_fft_64_stage_2_0_t338 * 32 +: 32] = FSM_fft_64_stage_2_0_t328 - FSM_fft_64_stage_2_0_t332;
    FSM_fft_64_stage_2_0_t340 = 32'b00000000000000000000000000001010 * 32'b00000000000000000000000000000100;
    FSM_fft_64_stage_2_0_t341 = FSM_fft_64_stage_2_0_t340[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t342 = FSM_fft_64_stage_2_0_t341[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t343 = FSM_fft_64_stage_2_0_t341[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t344 = FSM_fft_64_stage_2_0_t339[FSM_fft_64_stage_2_0_t343 * 32 +: 32];
    FSM_fft_64_stage_2_0_t345 = FSM_fft_64_stage_2_0_t341 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t346 = FSM_fft_64_stage_2_0_t345[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t347 = FSM_fft_64_stage_2_0_t346[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t348 = FSM_fft_64_stage_2_0_t339[FSM_fft_64_stage_2_0_t347 * 32 +: 32];
    FSM_fft_64_stage_2_0_t349 = FSM_fft_64_stage_2_0_t344 + FSM_fft_64_stage_2_0_t348;
    FSM_fft_64_stage_2_0_t350 = FSM_fft_64_stage_2_0_t349[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t351 = FSM_fft_64_stage_2_0_t339;
    FSM_fft_64_stage_2_0_t351[FSM_fft_64_stage_2_0_t342 * 32 +: 32] = FSM_fft_64_stage_2_0_t350;
    FSM_fft_64_stage_2_0_t352 = FSM_fft_64_stage_2_0_t341 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t353 = FSM_fft_64_stage_2_0_t352[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t354 = FSM_fft_64_stage_2_0_t353[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t355 = FSM_fft_64_stage_2_0_t351;
    FSM_fft_64_stage_2_0_t355[FSM_fft_64_stage_2_0_t354 * 32 +: 32] = FSM_fft_64_stage_2_0_t344 - FSM_fft_64_stage_2_0_t348;
    FSM_fft_64_stage_2_0_t356 = FSM_fft_64_stage_2_0_t341 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t357 = FSM_fft_64_stage_2_0_t356[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t358 = FSM_fft_64_stage_2_0_t357[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t359 = FSM_fft_64_stage_2_0_t341 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t360 = FSM_fft_64_stage_2_0_t359[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t361 = FSM_fft_64_stage_2_0_t360[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t362 = FSM_fft_64_stage_2_0_t339[FSM_fft_64_stage_2_0_t361 * 32 +: 32];
    FSM_fft_64_stage_2_0_t363 = FSM_fft_64_stage_2_0_t341 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t364 = FSM_fft_64_stage_2_0_t363[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t365 = FSM_fft_64_stage_2_0_t364[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t366 = FSM_fft_64_stage_2_0_t339[FSM_fft_64_stage_2_0_t365 * 32 +: 32];
    FSM_fft_64_stage_2_0_t367 = FSM_fft_64_stage_2_0_t362 + FSM_fft_64_stage_2_0_t366;
    FSM_fft_64_stage_2_0_t368 = FSM_fft_64_stage_2_0_t367[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t369 = FSM_fft_64_stage_2_0_t355;
    FSM_fft_64_stage_2_0_t369[FSM_fft_64_stage_2_0_t358 * 32 +: 32] = FSM_fft_64_stage_2_0_t368;
    FSM_fft_64_stage_2_0_t370 = FSM_fft_64_stage_2_0_t341 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t371 = FSM_fft_64_stage_2_0_t370[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t372 = FSM_fft_64_stage_2_0_t371[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t373 = FSM_fft_64_stage_2_0_t369;
    FSM_fft_64_stage_2_0_t373[FSM_fft_64_stage_2_0_t372 * 32 +: 32] = FSM_fft_64_stage_2_0_t362 - FSM_fft_64_stage_2_0_t366;
    FSM_fft_64_stage_2_0_t374 = 32'b00000000000000000000000000001011 * 32'b00000000000000000000000000000100;
    FSM_fft_64_stage_2_0_t375 = FSM_fft_64_stage_2_0_t374[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t376 = FSM_fft_64_stage_2_0_t375[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t377 = FSM_fft_64_stage_2_0_t375[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t378 = FSM_fft_64_stage_2_0_t373[FSM_fft_64_stage_2_0_t377 * 32 +: 32];
    FSM_fft_64_stage_2_0_t379 = FSM_fft_64_stage_2_0_t375 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t380 = FSM_fft_64_stage_2_0_t379[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t381 = FSM_fft_64_stage_2_0_t380[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t382 = FSM_fft_64_stage_2_0_t373[FSM_fft_64_stage_2_0_t381 * 32 +: 32];
    FSM_fft_64_stage_2_0_t383 = FSM_fft_64_stage_2_0_t378 + FSM_fft_64_stage_2_0_t382;
    FSM_fft_64_stage_2_0_t384 = FSM_fft_64_stage_2_0_t383[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t385 = FSM_fft_64_stage_2_0_t373;
    FSM_fft_64_stage_2_0_t385[FSM_fft_64_stage_2_0_t376 * 32 +: 32] = FSM_fft_64_stage_2_0_t384;
    FSM_fft_64_stage_2_0_t386 = FSM_fft_64_stage_2_0_t375 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t387 = FSM_fft_64_stage_2_0_t386[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t388 = FSM_fft_64_stage_2_0_t387[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t389 = FSM_fft_64_stage_2_0_t385;
    FSM_fft_64_stage_2_0_t389[FSM_fft_64_stage_2_0_t388 * 32 +: 32] = FSM_fft_64_stage_2_0_t378 - FSM_fft_64_stage_2_0_t382;
    FSM_fft_64_stage_2_0_t390 = FSM_fft_64_stage_2_0_t375 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t391 = FSM_fft_64_stage_2_0_t390[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t392 = FSM_fft_64_stage_2_0_t391[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t393 = FSM_fft_64_stage_2_0_t375 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t394 = FSM_fft_64_stage_2_0_t393[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t395 = FSM_fft_64_stage_2_0_t394[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t396 = FSM_fft_64_stage_2_0_t373[FSM_fft_64_stage_2_0_t395 * 32 +: 32];
    FSM_fft_64_stage_2_0_t397 = FSM_fft_64_stage_2_0_t375 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t398 = FSM_fft_64_stage_2_0_t397[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t399 = FSM_fft_64_stage_2_0_t398[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t400 = FSM_fft_64_stage_2_0_t373[FSM_fft_64_stage_2_0_t399 * 32 +: 32];
    FSM_fft_64_stage_2_0_t401 = FSM_fft_64_stage_2_0_t396 + FSM_fft_64_stage_2_0_t400;
    FSM_fft_64_stage_2_0_t402 = FSM_fft_64_stage_2_0_t401[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t403 = FSM_fft_64_stage_2_0_t389;
    FSM_fft_64_stage_2_0_t403[FSM_fft_64_stage_2_0_t392 * 32 +: 32] = FSM_fft_64_stage_2_0_t402;
    FSM_fft_64_stage_2_0_t404 = FSM_fft_64_stage_2_0_t375 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t405 = FSM_fft_64_stage_2_0_t404[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t406 = FSM_fft_64_stage_2_0_t405[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t407 = FSM_fft_64_stage_2_0_t403;
    FSM_fft_64_stage_2_0_t407[FSM_fft_64_stage_2_0_t406 * 32 +: 32] = FSM_fft_64_stage_2_0_t396 - FSM_fft_64_stage_2_0_t400;
    FSM_fft_64_stage_2_0_t408 = 32'b00000000000000000000000000001100 * 32'b00000000000000000000000000000100;
    FSM_fft_64_stage_2_0_t409 = FSM_fft_64_stage_2_0_t408[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t410 = FSM_fft_64_stage_2_0_t409[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t411 = FSM_fft_64_stage_2_0_t409[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t412 = FSM_fft_64_stage_2_0_t407[FSM_fft_64_stage_2_0_t411 * 32 +: 32];
    FSM_fft_64_stage_2_0_t413 = FSM_fft_64_stage_2_0_t409 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t414 = FSM_fft_64_stage_2_0_t413[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t415 = FSM_fft_64_stage_2_0_t414[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t416 = FSM_fft_64_stage_2_0_t407[FSM_fft_64_stage_2_0_t415 * 32 +: 32];
    FSM_fft_64_stage_2_0_t417 = FSM_fft_64_stage_2_0_t412 + FSM_fft_64_stage_2_0_t416;
    FSM_fft_64_stage_2_0_t418 = FSM_fft_64_stage_2_0_t417[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t419 = FSM_fft_64_stage_2_0_t407;
    FSM_fft_64_stage_2_0_t419[FSM_fft_64_stage_2_0_t410 * 32 +: 32] = FSM_fft_64_stage_2_0_t418;
    FSM_fft_64_stage_2_0_t420 = FSM_fft_64_stage_2_0_t409 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t421 = FSM_fft_64_stage_2_0_t420[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t422 = FSM_fft_64_stage_2_0_t421[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t423 = FSM_fft_64_stage_2_0_t419;
    FSM_fft_64_stage_2_0_t423[FSM_fft_64_stage_2_0_t422 * 32 +: 32] = FSM_fft_64_stage_2_0_t412 - FSM_fft_64_stage_2_0_t416;
    FSM_fft_64_stage_2_0_t424 = FSM_fft_64_stage_2_0_t409 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t425 = FSM_fft_64_stage_2_0_t424[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t426 = FSM_fft_64_stage_2_0_t425[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t427 = FSM_fft_64_stage_2_0_t409 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t428 = FSM_fft_64_stage_2_0_t427[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t429 = FSM_fft_64_stage_2_0_t428[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t430 = FSM_fft_64_stage_2_0_t407[FSM_fft_64_stage_2_0_t429 * 32 +: 32];
    FSM_fft_64_stage_2_0_t431 = FSM_fft_64_stage_2_0_t409 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t432 = FSM_fft_64_stage_2_0_t431[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t433 = FSM_fft_64_stage_2_0_t432[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t434 = FSM_fft_64_stage_2_0_t407[FSM_fft_64_stage_2_0_t433 * 32 +: 32];
    FSM_fft_64_stage_2_0_t435 = FSM_fft_64_stage_2_0_t430 + FSM_fft_64_stage_2_0_t434;
    FSM_fft_64_stage_2_0_t436 = FSM_fft_64_stage_2_0_t435[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t437 = FSM_fft_64_stage_2_0_t423;
    FSM_fft_64_stage_2_0_t437[FSM_fft_64_stage_2_0_t426 * 32 +: 32] = FSM_fft_64_stage_2_0_t436;
    FSM_fft_64_stage_2_0_t438 = FSM_fft_64_stage_2_0_t409 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t439 = FSM_fft_64_stage_2_0_t438[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t440 = FSM_fft_64_stage_2_0_t439[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t441 = FSM_fft_64_stage_2_0_t437;
    FSM_fft_64_stage_2_0_t441[FSM_fft_64_stage_2_0_t440 * 32 +: 32] = FSM_fft_64_stage_2_0_t430 - FSM_fft_64_stage_2_0_t434;
    FSM_fft_64_stage_2_0_t442 = 32'b00000000000000000000000000001101 * 32'b00000000000000000000000000000100;
    FSM_fft_64_stage_2_0_t443 = FSM_fft_64_stage_2_0_t442[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t444 = FSM_fft_64_stage_2_0_t443[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t445 = FSM_fft_64_stage_2_0_t443[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t446 = FSM_fft_64_stage_2_0_t441[FSM_fft_64_stage_2_0_t445 * 32 +: 32];
    FSM_fft_64_stage_2_0_t447 = FSM_fft_64_stage_2_0_t443 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t448 = FSM_fft_64_stage_2_0_t447[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t449 = FSM_fft_64_stage_2_0_t448[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t450 = FSM_fft_64_stage_2_0_t441[FSM_fft_64_stage_2_0_t449 * 32 +: 32];
    FSM_fft_64_stage_2_0_t451 = FSM_fft_64_stage_2_0_t446 + FSM_fft_64_stage_2_0_t450;
    FSM_fft_64_stage_2_0_t452 = FSM_fft_64_stage_2_0_t451[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t453 = FSM_fft_64_stage_2_0_t441;
    FSM_fft_64_stage_2_0_t453[FSM_fft_64_stage_2_0_t444 * 32 +: 32] = FSM_fft_64_stage_2_0_t452;
    FSM_fft_64_stage_2_0_t454 = FSM_fft_64_stage_2_0_t443 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t455 = FSM_fft_64_stage_2_0_t454[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t456 = FSM_fft_64_stage_2_0_t455[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t457 = FSM_fft_64_stage_2_0_t453;
    FSM_fft_64_stage_2_0_t457[FSM_fft_64_stage_2_0_t456 * 32 +: 32] = FSM_fft_64_stage_2_0_t446 - FSM_fft_64_stage_2_0_t450;
    FSM_fft_64_stage_2_0_t458 = FSM_fft_64_stage_2_0_t443 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t459 = FSM_fft_64_stage_2_0_t458[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t460 = FSM_fft_64_stage_2_0_t459[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t461 = FSM_fft_64_stage_2_0_t443 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t462 = FSM_fft_64_stage_2_0_t461[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t463 = FSM_fft_64_stage_2_0_t462[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t464 = FSM_fft_64_stage_2_0_t441[FSM_fft_64_stage_2_0_t463 * 32 +: 32];
    FSM_fft_64_stage_2_0_t465 = FSM_fft_64_stage_2_0_t443 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t466 = FSM_fft_64_stage_2_0_t465[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t467 = FSM_fft_64_stage_2_0_t466[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t468 = FSM_fft_64_stage_2_0_t441[FSM_fft_64_stage_2_0_t467 * 32 +: 32];
    FSM_fft_64_stage_2_0_t469 = FSM_fft_64_stage_2_0_t464 + FSM_fft_64_stage_2_0_t468;
    FSM_fft_64_stage_2_0_t470 = FSM_fft_64_stage_2_0_t469[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t471 = FSM_fft_64_stage_2_0_t457;
    FSM_fft_64_stage_2_0_t471[FSM_fft_64_stage_2_0_t460 * 32 +: 32] = FSM_fft_64_stage_2_0_t470;
    FSM_fft_64_stage_2_0_t472 = FSM_fft_64_stage_2_0_t443 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t473 = FSM_fft_64_stage_2_0_t472[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t474 = FSM_fft_64_stage_2_0_t473[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t475 = FSM_fft_64_stage_2_0_t471;
    FSM_fft_64_stage_2_0_t475[FSM_fft_64_stage_2_0_t474 * 32 +: 32] = FSM_fft_64_stage_2_0_t464 - FSM_fft_64_stage_2_0_t468;
    FSM_fft_64_stage_2_0_t476 = 32'b00000000000000000000000000001110 * 32'b00000000000000000000000000000100;
    FSM_fft_64_stage_2_0_t477 = FSM_fft_64_stage_2_0_t476[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t478 = FSM_fft_64_stage_2_0_t477[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t479 = FSM_fft_64_stage_2_0_t477[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t480 = FSM_fft_64_stage_2_0_t475[FSM_fft_64_stage_2_0_t479 * 32 +: 32];
    FSM_fft_64_stage_2_0_t481 = FSM_fft_64_stage_2_0_t477 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t482 = FSM_fft_64_stage_2_0_t481[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t483 = FSM_fft_64_stage_2_0_t482[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t484 = FSM_fft_64_stage_2_0_t475[FSM_fft_64_stage_2_0_t483 * 32 +: 32];
    FSM_fft_64_stage_2_0_t485 = FSM_fft_64_stage_2_0_t480 + FSM_fft_64_stage_2_0_t484;
    FSM_fft_64_stage_2_0_t486 = FSM_fft_64_stage_2_0_t485[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t487 = FSM_fft_64_stage_2_0_t475;
    FSM_fft_64_stage_2_0_t487[FSM_fft_64_stage_2_0_t478 * 32 +: 32] = FSM_fft_64_stage_2_0_t486;
    FSM_fft_64_stage_2_0_t488 = FSM_fft_64_stage_2_0_t477 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t489 = FSM_fft_64_stage_2_0_t488[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t490 = FSM_fft_64_stage_2_0_t489[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t491 = FSM_fft_64_stage_2_0_t487;
    FSM_fft_64_stage_2_0_t491[FSM_fft_64_stage_2_0_t490 * 32 +: 32] = FSM_fft_64_stage_2_0_t480 - FSM_fft_64_stage_2_0_t484;
    FSM_fft_64_stage_2_0_t492 = FSM_fft_64_stage_2_0_t477 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t493 = FSM_fft_64_stage_2_0_t492[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t494 = FSM_fft_64_stage_2_0_t493[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t495 = FSM_fft_64_stage_2_0_t477 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t496 = FSM_fft_64_stage_2_0_t495[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t497 = FSM_fft_64_stage_2_0_t496[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t498 = FSM_fft_64_stage_2_0_t475[FSM_fft_64_stage_2_0_t497 * 32 +: 32];
    FSM_fft_64_stage_2_0_t499 = FSM_fft_64_stage_2_0_t477 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t500 = FSM_fft_64_stage_2_0_t499[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t501 = FSM_fft_64_stage_2_0_t500[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t502 = FSM_fft_64_stage_2_0_t475[FSM_fft_64_stage_2_0_t501 * 32 +: 32];
    FSM_fft_64_stage_2_0_t503 = FSM_fft_64_stage_2_0_t498 + FSM_fft_64_stage_2_0_t502;
    FSM_fft_64_stage_2_0_t504 = FSM_fft_64_stage_2_0_t503[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t505 = FSM_fft_64_stage_2_0_t491;
    FSM_fft_64_stage_2_0_t505[FSM_fft_64_stage_2_0_t494 * 32 +: 32] = FSM_fft_64_stage_2_0_t504;
    FSM_fft_64_stage_2_0_t506 = FSM_fft_64_stage_2_0_t477 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t507 = FSM_fft_64_stage_2_0_t506[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t508 = FSM_fft_64_stage_2_0_t507[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t509 = FSM_fft_64_stage_2_0_t505;
    FSM_fft_64_stage_2_0_t509[FSM_fft_64_stage_2_0_t508 * 32 +: 32] = FSM_fft_64_stage_2_0_t498 - FSM_fft_64_stage_2_0_t502;
    FSM_fft_64_stage_2_0_t510 = 32'b00000000000000000000000000001111 * 32'b00000000000000000000000000000100;
    FSM_fft_64_stage_2_0_t511 = FSM_fft_64_stage_2_0_t510[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t512 = FSM_fft_64_stage_2_0_t511[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t513 = FSM_fft_64_stage_2_0_t511[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t514 = FSM_fft_64_stage_2_0_t509[FSM_fft_64_stage_2_0_t513 * 32 +: 32];
    FSM_fft_64_stage_2_0_t515 = FSM_fft_64_stage_2_0_t511 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t516 = FSM_fft_64_stage_2_0_t515[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t517 = FSM_fft_64_stage_2_0_t516[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t518 = FSM_fft_64_stage_2_0_t509[FSM_fft_64_stage_2_0_t517 * 32 +: 32];
    FSM_fft_64_stage_2_0_t519 = FSM_fft_64_stage_2_0_t514 + FSM_fft_64_stage_2_0_t518;
    FSM_fft_64_stage_2_0_t520 = FSM_fft_64_stage_2_0_t519[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t521 = FSM_fft_64_stage_2_0_t509;
    FSM_fft_64_stage_2_0_t521[FSM_fft_64_stage_2_0_t512 * 32 +: 32] = FSM_fft_64_stage_2_0_t520;
    FSM_fft_64_stage_2_0_t522 = FSM_fft_64_stage_2_0_t511 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t523 = FSM_fft_64_stage_2_0_t522[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t524 = FSM_fft_64_stage_2_0_t523[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t525 = FSM_fft_64_stage_2_0_t521;
    FSM_fft_64_stage_2_0_t525[FSM_fft_64_stage_2_0_t524 * 32 +: 32] = FSM_fft_64_stage_2_0_t514 - FSM_fft_64_stage_2_0_t518;
    FSM_fft_64_stage_2_0_t526 = FSM_fft_64_stage_2_0_t511 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t527 = FSM_fft_64_stage_2_0_t526[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t528 = FSM_fft_64_stage_2_0_t527[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t529 = FSM_fft_64_stage_2_0_t511 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t530 = FSM_fft_64_stage_2_0_t529[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t531 = FSM_fft_64_stage_2_0_t530[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t532 = FSM_fft_64_stage_2_0_t509[FSM_fft_64_stage_2_0_t531 * 32 +: 32];
    FSM_fft_64_stage_2_0_t533 = FSM_fft_64_stage_2_0_t511 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t534 = FSM_fft_64_stage_2_0_t533[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t535 = FSM_fft_64_stage_2_0_t534[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t536 = FSM_fft_64_stage_2_0_t509[FSM_fft_64_stage_2_0_t535 * 32 +: 32];
    FSM_fft_64_stage_2_0_t537 = FSM_fft_64_stage_2_0_t532 + FSM_fft_64_stage_2_0_t536;
    FSM_fft_64_stage_2_0_t538 = FSM_fft_64_stage_2_0_t537[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t539 = FSM_fft_64_stage_2_0_t525;
    FSM_fft_64_stage_2_0_t539[FSM_fft_64_stage_2_0_t528 * 32 +: 32] = FSM_fft_64_stage_2_0_t538;
    FSM_fft_64_stage_2_0_t540 = FSM_fft_64_stage_2_0_t511 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t541 = FSM_fft_64_stage_2_0_t540[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t542 = FSM_fft_64_stage_2_0_t541[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t543 = FSM_fft_64_stage_2_0_t539;
    FSM_fft_64_stage_2_0_t543[FSM_fft_64_stage_2_0_t542 * 32 +: 32] = FSM_fft_64_stage_2_0_t532 - FSM_fft_64_stage_2_0_t536;
    FSM_fft_64_stage_2_0_t544 = FSM_fft_64_stage_2_0_t1[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t545 = FSM_fft_64_stage_2_0_t1[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t546 = i_data_in_imag[FSM_fft_64_stage_2_0_t545 * 32 +: 32];
    FSM_fft_64_stage_2_0_t547 = FSM_fft_64_stage_2_0_t1 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t548 = FSM_fft_64_stage_2_0_t547[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t549 = FSM_fft_64_stage_2_0_t548[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t550 = i_data_in_imag[FSM_fft_64_stage_2_0_t549 * 32 +: 32];
    FSM_fft_64_stage_2_0_t551 = FSM_fft_64_stage_2_0_t546 + FSM_fft_64_stage_2_0_t550;
    FSM_fft_64_stage_2_0_t552 = FSM_fft_64_stage_2_0_t551[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t553 = i_data_in_imag;
    FSM_fft_64_stage_2_0_t553[FSM_fft_64_stage_2_0_t544 * 32 +: 32] = FSM_fft_64_stage_2_0_t552;
    FSM_fft_64_stage_2_0_t554 = FSM_fft_64_stage_2_0_t1 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t555 = FSM_fft_64_stage_2_0_t554[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t556 = FSM_fft_64_stage_2_0_t555[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t557 = FSM_fft_64_stage_2_0_t553;
    FSM_fft_64_stage_2_0_t557[FSM_fft_64_stage_2_0_t556 * 32 +: 32] = FSM_fft_64_stage_2_0_t546 - FSM_fft_64_stage_2_0_t550;
    FSM_fft_64_stage_2_0_t558 = FSM_fft_64_stage_2_0_t1 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t559 = FSM_fft_64_stage_2_0_t558[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t560 = FSM_fft_64_stage_2_0_t559[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t561 = FSM_fft_64_stage_2_0_t1 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t562 = FSM_fft_64_stage_2_0_t561[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t563 = FSM_fft_64_stage_2_0_t562[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t564 = i_data_in_imag[FSM_fft_64_stage_2_0_t563 * 32 +: 32];
    FSM_fft_64_stage_2_0_t565 = FSM_fft_64_stage_2_0_t1 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t566 = FSM_fft_64_stage_2_0_t565[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t567 = FSM_fft_64_stage_2_0_t566[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t568 = i_data_in_imag[FSM_fft_64_stage_2_0_t567 * 32 +: 32];
    FSM_fft_64_stage_2_0_t569 = FSM_fft_64_stage_2_0_t564 + FSM_fft_64_stage_2_0_t568;
    FSM_fft_64_stage_2_0_t570 = FSM_fft_64_stage_2_0_t569[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t571 = FSM_fft_64_stage_2_0_t557;
    FSM_fft_64_stage_2_0_t571[FSM_fft_64_stage_2_0_t560 * 32 +: 32] = FSM_fft_64_stage_2_0_t570;
    FSM_fft_64_stage_2_0_t572 = FSM_fft_64_stage_2_0_t1 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t573 = FSM_fft_64_stage_2_0_t572[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t574 = FSM_fft_64_stage_2_0_t573[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t575 = FSM_fft_64_stage_2_0_t571;
    FSM_fft_64_stage_2_0_t575[FSM_fft_64_stage_2_0_t574 * 32 +: 32] = FSM_fft_64_stage_2_0_t564 - FSM_fft_64_stage_2_0_t568;
    FSM_fft_64_stage_2_0_t576 = FSM_fft_64_stage_2_0_t35[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t577 = FSM_fft_64_stage_2_0_t35[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t578 = FSM_fft_64_stage_2_0_t575[FSM_fft_64_stage_2_0_t577 * 32 +: 32];
    FSM_fft_64_stage_2_0_t579 = FSM_fft_64_stage_2_0_t35 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t580 = FSM_fft_64_stage_2_0_t579[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t581 = FSM_fft_64_stage_2_0_t580[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t582 = FSM_fft_64_stage_2_0_t575[FSM_fft_64_stage_2_0_t581 * 32 +: 32];
    FSM_fft_64_stage_2_0_t583 = FSM_fft_64_stage_2_0_t578 + FSM_fft_64_stage_2_0_t582;
    FSM_fft_64_stage_2_0_t584 = FSM_fft_64_stage_2_0_t583[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t585 = FSM_fft_64_stage_2_0_t575;
    FSM_fft_64_stage_2_0_t585[FSM_fft_64_stage_2_0_t576 * 32 +: 32] = FSM_fft_64_stage_2_0_t584;
    FSM_fft_64_stage_2_0_t586 = FSM_fft_64_stage_2_0_t35 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t587 = FSM_fft_64_stage_2_0_t586[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t588 = FSM_fft_64_stage_2_0_t587[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t589 = FSM_fft_64_stage_2_0_t585;
    FSM_fft_64_stage_2_0_t589[FSM_fft_64_stage_2_0_t588 * 32 +: 32] = FSM_fft_64_stage_2_0_t578 - FSM_fft_64_stage_2_0_t582;
    FSM_fft_64_stage_2_0_t590 = FSM_fft_64_stage_2_0_t35 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t591 = FSM_fft_64_stage_2_0_t590[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t592 = FSM_fft_64_stage_2_0_t591[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t593 = FSM_fft_64_stage_2_0_t35 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t594 = FSM_fft_64_stage_2_0_t593[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t595 = FSM_fft_64_stage_2_0_t594[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t596 = FSM_fft_64_stage_2_0_t575[FSM_fft_64_stage_2_0_t595 * 32 +: 32];
    FSM_fft_64_stage_2_0_t597 = FSM_fft_64_stage_2_0_t35 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t598 = FSM_fft_64_stage_2_0_t597[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t599 = FSM_fft_64_stage_2_0_t598[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t600 = FSM_fft_64_stage_2_0_t575[FSM_fft_64_stage_2_0_t599 * 32 +: 32];
    FSM_fft_64_stage_2_0_t601 = FSM_fft_64_stage_2_0_t596 + FSM_fft_64_stage_2_0_t600;
    FSM_fft_64_stage_2_0_t602 = FSM_fft_64_stage_2_0_t601[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t603 = FSM_fft_64_stage_2_0_t589;
    FSM_fft_64_stage_2_0_t603[FSM_fft_64_stage_2_0_t592 * 32 +: 32] = FSM_fft_64_stage_2_0_t602;
    FSM_fft_64_stage_2_0_t604 = FSM_fft_64_stage_2_0_t35 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t605 = FSM_fft_64_stage_2_0_t604[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t606 = FSM_fft_64_stage_2_0_t605[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t607 = FSM_fft_64_stage_2_0_t603;
    FSM_fft_64_stage_2_0_t607[FSM_fft_64_stage_2_0_t606 * 32 +: 32] = FSM_fft_64_stage_2_0_t596 - FSM_fft_64_stage_2_0_t600;
    FSM_fft_64_stage_2_0_t608 = FSM_fft_64_stage_2_0_t69[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t609 = FSM_fft_64_stage_2_0_t69[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t610 = FSM_fft_64_stage_2_0_t607[FSM_fft_64_stage_2_0_t609 * 32 +: 32];
    FSM_fft_64_stage_2_0_t611 = FSM_fft_64_stage_2_0_t69 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t612 = FSM_fft_64_stage_2_0_t611[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t613 = FSM_fft_64_stage_2_0_t612[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t614 = FSM_fft_64_stage_2_0_t607[FSM_fft_64_stage_2_0_t613 * 32 +: 32];
    FSM_fft_64_stage_2_0_t615 = FSM_fft_64_stage_2_0_t610 + FSM_fft_64_stage_2_0_t614;
    FSM_fft_64_stage_2_0_t616 = FSM_fft_64_stage_2_0_t615[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t617 = FSM_fft_64_stage_2_0_t607;
    FSM_fft_64_stage_2_0_t617[FSM_fft_64_stage_2_0_t608 * 32 +: 32] = FSM_fft_64_stage_2_0_t616;
    FSM_fft_64_stage_2_0_t618 = FSM_fft_64_stage_2_0_t69 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t619 = FSM_fft_64_stage_2_0_t618[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t620 = FSM_fft_64_stage_2_0_t619[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t621 = FSM_fft_64_stage_2_0_t617;
    FSM_fft_64_stage_2_0_t621[FSM_fft_64_stage_2_0_t620 * 32 +: 32] = FSM_fft_64_stage_2_0_t610 - FSM_fft_64_stage_2_0_t614;
    FSM_fft_64_stage_2_0_t622 = FSM_fft_64_stage_2_0_t69 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t623 = FSM_fft_64_stage_2_0_t622[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t624 = FSM_fft_64_stage_2_0_t623[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t625 = FSM_fft_64_stage_2_0_t69 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t626 = FSM_fft_64_stage_2_0_t625[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t627 = FSM_fft_64_stage_2_0_t626[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t628 = FSM_fft_64_stage_2_0_t607[FSM_fft_64_stage_2_0_t627 * 32 +: 32];
    FSM_fft_64_stage_2_0_t629 = FSM_fft_64_stage_2_0_t69 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t630 = FSM_fft_64_stage_2_0_t629[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t631 = FSM_fft_64_stage_2_0_t630[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t632 = FSM_fft_64_stage_2_0_t607[FSM_fft_64_stage_2_0_t631 * 32 +: 32];
    FSM_fft_64_stage_2_0_t633 = FSM_fft_64_stage_2_0_t628 + FSM_fft_64_stage_2_0_t632;
    FSM_fft_64_stage_2_0_t634 = FSM_fft_64_stage_2_0_t633[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t635 = FSM_fft_64_stage_2_0_t621;
    FSM_fft_64_stage_2_0_t635[FSM_fft_64_stage_2_0_t624 * 32 +: 32] = FSM_fft_64_stage_2_0_t634;
    FSM_fft_64_stage_2_0_t636 = FSM_fft_64_stage_2_0_t69 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t637 = FSM_fft_64_stage_2_0_t636[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t638 = FSM_fft_64_stage_2_0_t637[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t639 = FSM_fft_64_stage_2_0_t635;
    FSM_fft_64_stage_2_0_t639[FSM_fft_64_stage_2_0_t638 * 32 +: 32] = FSM_fft_64_stage_2_0_t628 - FSM_fft_64_stage_2_0_t632;
    FSM_fft_64_stage_2_0_t640 = FSM_fft_64_stage_2_0_t103[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t641 = FSM_fft_64_stage_2_0_t103[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t642 = FSM_fft_64_stage_2_0_t639[FSM_fft_64_stage_2_0_t641 * 32 +: 32];
    FSM_fft_64_stage_2_0_t643 = FSM_fft_64_stage_2_0_t103 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t644 = FSM_fft_64_stage_2_0_t643[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t645 = FSM_fft_64_stage_2_0_t644[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t646 = FSM_fft_64_stage_2_0_t639[FSM_fft_64_stage_2_0_t645 * 32 +: 32];
    FSM_fft_64_stage_2_0_t647 = FSM_fft_64_stage_2_0_t642 + FSM_fft_64_stage_2_0_t646;
    FSM_fft_64_stage_2_0_t648 = FSM_fft_64_stage_2_0_t647[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t649 = FSM_fft_64_stage_2_0_t639;
    FSM_fft_64_stage_2_0_t649[FSM_fft_64_stage_2_0_t640 * 32 +: 32] = FSM_fft_64_stage_2_0_t648;
    FSM_fft_64_stage_2_0_t650 = FSM_fft_64_stage_2_0_t103 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t651 = FSM_fft_64_stage_2_0_t650[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t652 = FSM_fft_64_stage_2_0_t651[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t653 = FSM_fft_64_stage_2_0_t649;
    FSM_fft_64_stage_2_0_t653[FSM_fft_64_stage_2_0_t652 * 32 +: 32] = FSM_fft_64_stage_2_0_t642 - FSM_fft_64_stage_2_0_t646;
    FSM_fft_64_stage_2_0_t654 = FSM_fft_64_stage_2_0_t103 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t655 = FSM_fft_64_stage_2_0_t654[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t656 = FSM_fft_64_stage_2_0_t655[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t657 = FSM_fft_64_stage_2_0_t103 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t658 = FSM_fft_64_stage_2_0_t657[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t659 = FSM_fft_64_stage_2_0_t658[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t660 = FSM_fft_64_stage_2_0_t639[FSM_fft_64_stage_2_0_t659 * 32 +: 32];
    FSM_fft_64_stage_2_0_t661 = FSM_fft_64_stage_2_0_t103 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t662 = FSM_fft_64_stage_2_0_t661[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t663 = FSM_fft_64_stage_2_0_t662[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t664 = FSM_fft_64_stage_2_0_t639[FSM_fft_64_stage_2_0_t663 * 32 +: 32];
    FSM_fft_64_stage_2_0_t665 = FSM_fft_64_stage_2_0_t660 + FSM_fft_64_stage_2_0_t664;
    FSM_fft_64_stage_2_0_t666 = FSM_fft_64_stage_2_0_t665[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t667 = FSM_fft_64_stage_2_0_t653;
    FSM_fft_64_stage_2_0_t667[FSM_fft_64_stage_2_0_t656 * 32 +: 32] = FSM_fft_64_stage_2_0_t666;
    FSM_fft_64_stage_2_0_t668 = FSM_fft_64_stage_2_0_t103 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t669 = FSM_fft_64_stage_2_0_t668[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t670 = FSM_fft_64_stage_2_0_t669[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t671 = FSM_fft_64_stage_2_0_t667;
    FSM_fft_64_stage_2_0_t671[FSM_fft_64_stage_2_0_t670 * 32 +: 32] = FSM_fft_64_stage_2_0_t660 - FSM_fft_64_stage_2_0_t664;
    FSM_fft_64_stage_2_0_t672 = FSM_fft_64_stage_2_0_t137[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t673 = FSM_fft_64_stage_2_0_t137[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t674 = FSM_fft_64_stage_2_0_t671[FSM_fft_64_stage_2_0_t673 * 32 +: 32];
    FSM_fft_64_stage_2_0_t675 = FSM_fft_64_stage_2_0_t137 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t676 = FSM_fft_64_stage_2_0_t675[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t677 = FSM_fft_64_stage_2_0_t676[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t678 = FSM_fft_64_stage_2_0_t671[FSM_fft_64_stage_2_0_t677 * 32 +: 32];
    FSM_fft_64_stage_2_0_t679 = FSM_fft_64_stage_2_0_t674 + FSM_fft_64_stage_2_0_t678;
    FSM_fft_64_stage_2_0_t680 = FSM_fft_64_stage_2_0_t679[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t681 = FSM_fft_64_stage_2_0_t671;
    FSM_fft_64_stage_2_0_t681[FSM_fft_64_stage_2_0_t672 * 32 +: 32] = FSM_fft_64_stage_2_0_t680;
    FSM_fft_64_stage_2_0_t682 = FSM_fft_64_stage_2_0_t137 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t683 = FSM_fft_64_stage_2_0_t682[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t684 = FSM_fft_64_stage_2_0_t683[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t685 = FSM_fft_64_stage_2_0_t681;
    FSM_fft_64_stage_2_0_t685[FSM_fft_64_stage_2_0_t684 * 32 +: 32] = FSM_fft_64_stage_2_0_t674 - FSM_fft_64_stage_2_0_t678;
    FSM_fft_64_stage_2_0_t686 = FSM_fft_64_stage_2_0_t137 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t687 = FSM_fft_64_stage_2_0_t686[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t688 = FSM_fft_64_stage_2_0_t687[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t689 = FSM_fft_64_stage_2_0_t137 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t690 = FSM_fft_64_stage_2_0_t689[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t691 = FSM_fft_64_stage_2_0_t690[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t692 = FSM_fft_64_stage_2_0_t671[FSM_fft_64_stage_2_0_t691 * 32 +: 32];
    FSM_fft_64_stage_2_0_t693 = FSM_fft_64_stage_2_0_t137 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t694 = FSM_fft_64_stage_2_0_t693[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t695 = FSM_fft_64_stage_2_0_t694[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t696 = FSM_fft_64_stage_2_0_t671[FSM_fft_64_stage_2_0_t695 * 32 +: 32];
    FSM_fft_64_stage_2_0_t697 = FSM_fft_64_stage_2_0_t692 + FSM_fft_64_stage_2_0_t696;
    FSM_fft_64_stage_2_0_t698 = FSM_fft_64_stage_2_0_t697[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t699 = FSM_fft_64_stage_2_0_t685;
    FSM_fft_64_stage_2_0_t699[FSM_fft_64_stage_2_0_t688 * 32 +: 32] = FSM_fft_64_stage_2_0_t698;
    FSM_fft_64_stage_2_0_t700 = FSM_fft_64_stage_2_0_t137 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t701 = FSM_fft_64_stage_2_0_t700[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t702 = FSM_fft_64_stage_2_0_t701[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t703 = FSM_fft_64_stage_2_0_t699;
    FSM_fft_64_stage_2_0_t703[FSM_fft_64_stage_2_0_t702 * 32 +: 32] = FSM_fft_64_stage_2_0_t692 - FSM_fft_64_stage_2_0_t696;
    FSM_fft_64_stage_2_0_t704 = FSM_fft_64_stage_2_0_t171[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t705 = FSM_fft_64_stage_2_0_t171[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t706 = FSM_fft_64_stage_2_0_t703[FSM_fft_64_stage_2_0_t705 * 32 +: 32];
    FSM_fft_64_stage_2_0_t707 = FSM_fft_64_stage_2_0_t171 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t708 = FSM_fft_64_stage_2_0_t707[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t709 = FSM_fft_64_stage_2_0_t708[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t710 = FSM_fft_64_stage_2_0_t703[FSM_fft_64_stage_2_0_t709 * 32 +: 32];
    FSM_fft_64_stage_2_0_t711 = FSM_fft_64_stage_2_0_t706 + FSM_fft_64_stage_2_0_t710;
    FSM_fft_64_stage_2_0_t712 = FSM_fft_64_stage_2_0_t711[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t713 = FSM_fft_64_stage_2_0_t703;
    FSM_fft_64_stage_2_0_t713[FSM_fft_64_stage_2_0_t704 * 32 +: 32] = FSM_fft_64_stage_2_0_t712;
    FSM_fft_64_stage_2_0_t714 = FSM_fft_64_stage_2_0_t171 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t715 = FSM_fft_64_stage_2_0_t714[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t716 = FSM_fft_64_stage_2_0_t715[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t717 = FSM_fft_64_stage_2_0_t713;
    FSM_fft_64_stage_2_0_t717[FSM_fft_64_stage_2_0_t716 * 32 +: 32] = FSM_fft_64_stage_2_0_t706 - FSM_fft_64_stage_2_0_t710;
    FSM_fft_64_stage_2_0_t718 = FSM_fft_64_stage_2_0_t171 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t719 = FSM_fft_64_stage_2_0_t718[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t720 = FSM_fft_64_stage_2_0_t719[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t721 = FSM_fft_64_stage_2_0_t171 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t722 = FSM_fft_64_stage_2_0_t721[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t723 = FSM_fft_64_stage_2_0_t722[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t724 = FSM_fft_64_stage_2_0_t703[FSM_fft_64_stage_2_0_t723 * 32 +: 32];
    FSM_fft_64_stage_2_0_t725 = FSM_fft_64_stage_2_0_t171 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t726 = FSM_fft_64_stage_2_0_t725[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t727 = FSM_fft_64_stage_2_0_t726[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t728 = FSM_fft_64_stage_2_0_t703[FSM_fft_64_stage_2_0_t727 * 32 +: 32];
    FSM_fft_64_stage_2_0_t729 = FSM_fft_64_stage_2_0_t724 + FSM_fft_64_stage_2_0_t728;
    FSM_fft_64_stage_2_0_t730 = FSM_fft_64_stage_2_0_t729[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t731 = FSM_fft_64_stage_2_0_t717;
    FSM_fft_64_stage_2_0_t731[FSM_fft_64_stage_2_0_t720 * 32 +: 32] = FSM_fft_64_stage_2_0_t730;
    FSM_fft_64_stage_2_0_t732 = FSM_fft_64_stage_2_0_t171 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t733 = FSM_fft_64_stage_2_0_t732[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t734 = FSM_fft_64_stage_2_0_t733[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t735 = FSM_fft_64_stage_2_0_t731;
    FSM_fft_64_stage_2_0_t735[FSM_fft_64_stage_2_0_t734 * 32 +: 32] = FSM_fft_64_stage_2_0_t724 - FSM_fft_64_stage_2_0_t728;
    FSM_fft_64_stage_2_0_t736 = FSM_fft_64_stage_2_0_t205[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t737 = FSM_fft_64_stage_2_0_t205[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t738 = FSM_fft_64_stage_2_0_t735[FSM_fft_64_stage_2_0_t737 * 32 +: 32];
    FSM_fft_64_stage_2_0_t739 = FSM_fft_64_stage_2_0_t205 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t740 = FSM_fft_64_stage_2_0_t739[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t741 = FSM_fft_64_stage_2_0_t740[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t742 = FSM_fft_64_stage_2_0_t735[FSM_fft_64_stage_2_0_t741 * 32 +: 32];
    FSM_fft_64_stage_2_0_t743 = FSM_fft_64_stage_2_0_t738 + FSM_fft_64_stage_2_0_t742;
    FSM_fft_64_stage_2_0_t744 = FSM_fft_64_stage_2_0_t743[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t745 = FSM_fft_64_stage_2_0_t735;
    FSM_fft_64_stage_2_0_t745[FSM_fft_64_stage_2_0_t736 * 32 +: 32] = FSM_fft_64_stage_2_0_t744;
    FSM_fft_64_stage_2_0_t746 = FSM_fft_64_stage_2_0_t205 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t747 = FSM_fft_64_stage_2_0_t746[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t748 = FSM_fft_64_stage_2_0_t747[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t749 = FSM_fft_64_stage_2_0_t745;
    FSM_fft_64_stage_2_0_t749[FSM_fft_64_stage_2_0_t748 * 32 +: 32] = FSM_fft_64_stage_2_0_t738 - FSM_fft_64_stage_2_0_t742;
    FSM_fft_64_stage_2_0_t750 = FSM_fft_64_stage_2_0_t205 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t751 = FSM_fft_64_stage_2_0_t750[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t752 = FSM_fft_64_stage_2_0_t751[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t753 = FSM_fft_64_stage_2_0_t205 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t754 = FSM_fft_64_stage_2_0_t753[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t755 = FSM_fft_64_stage_2_0_t754[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t756 = FSM_fft_64_stage_2_0_t735[FSM_fft_64_stage_2_0_t755 * 32 +: 32];
    FSM_fft_64_stage_2_0_t757 = FSM_fft_64_stage_2_0_t205 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t758 = FSM_fft_64_stage_2_0_t757[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t759 = FSM_fft_64_stage_2_0_t758[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t760 = FSM_fft_64_stage_2_0_t735[FSM_fft_64_stage_2_0_t759 * 32 +: 32];
    FSM_fft_64_stage_2_0_t761 = FSM_fft_64_stage_2_0_t756 + FSM_fft_64_stage_2_0_t760;
    FSM_fft_64_stage_2_0_t762 = FSM_fft_64_stage_2_0_t761[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t763 = FSM_fft_64_stage_2_0_t749;
    FSM_fft_64_stage_2_0_t763[FSM_fft_64_stage_2_0_t752 * 32 +: 32] = FSM_fft_64_stage_2_0_t762;
    FSM_fft_64_stage_2_0_t764 = FSM_fft_64_stage_2_0_t205 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t765 = FSM_fft_64_stage_2_0_t764[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t766 = FSM_fft_64_stage_2_0_t765[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t767 = FSM_fft_64_stage_2_0_t763;
    FSM_fft_64_stage_2_0_t767[FSM_fft_64_stage_2_0_t766 * 32 +: 32] = FSM_fft_64_stage_2_0_t756 - FSM_fft_64_stage_2_0_t760;
    FSM_fft_64_stage_2_0_t768 = FSM_fft_64_stage_2_0_t239[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t769 = FSM_fft_64_stage_2_0_t239[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t770 = FSM_fft_64_stage_2_0_t767[FSM_fft_64_stage_2_0_t769 * 32 +: 32];
    FSM_fft_64_stage_2_0_t771 = FSM_fft_64_stage_2_0_t239 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t772 = FSM_fft_64_stage_2_0_t771[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t773 = FSM_fft_64_stage_2_0_t772[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t774 = FSM_fft_64_stage_2_0_t767[FSM_fft_64_stage_2_0_t773 * 32 +: 32];
    FSM_fft_64_stage_2_0_t775 = FSM_fft_64_stage_2_0_t770 + FSM_fft_64_stage_2_0_t774;
    FSM_fft_64_stage_2_0_t776 = FSM_fft_64_stage_2_0_t775[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t777 = FSM_fft_64_stage_2_0_t767;
    FSM_fft_64_stage_2_0_t777[FSM_fft_64_stage_2_0_t768 * 32 +: 32] = FSM_fft_64_stage_2_0_t776;
    FSM_fft_64_stage_2_0_t778 = FSM_fft_64_stage_2_0_t239 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t779 = FSM_fft_64_stage_2_0_t778[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t780 = FSM_fft_64_stage_2_0_t779[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t781 = FSM_fft_64_stage_2_0_t777;
    FSM_fft_64_stage_2_0_t781[FSM_fft_64_stage_2_0_t780 * 32 +: 32] = FSM_fft_64_stage_2_0_t770 - FSM_fft_64_stage_2_0_t774;
    FSM_fft_64_stage_2_0_t782 = FSM_fft_64_stage_2_0_t239 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t783 = FSM_fft_64_stage_2_0_t782[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t784 = FSM_fft_64_stage_2_0_t783[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t785 = FSM_fft_64_stage_2_0_t239 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t786 = FSM_fft_64_stage_2_0_t785[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t787 = FSM_fft_64_stage_2_0_t786[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t788 = FSM_fft_64_stage_2_0_t767[FSM_fft_64_stage_2_0_t787 * 32 +: 32];
    FSM_fft_64_stage_2_0_t789 = FSM_fft_64_stage_2_0_t239 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t790 = FSM_fft_64_stage_2_0_t789[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t791 = FSM_fft_64_stage_2_0_t790[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t792 = FSM_fft_64_stage_2_0_t767[FSM_fft_64_stage_2_0_t791 * 32 +: 32];
    FSM_fft_64_stage_2_0_t793 = FSM_fft_64_stage_2_0_t788 + FSM_fft_64_stage_2_0_t792;
    FSM_fft_64_stage_2_0_t794 = FSM_fft_64_stage_2_0_t793[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t795 = FSM_fft_64_stage_2_0_t781;
    FSM_fft_64_stage_2_0_t795[FSM_fft_64_stage_2_0_t784 * 32 +: 32] = FSM_fft_64_stage_2_0_t794;
    FSM_fft_64_stage_2_0_t796 = FSM_fft_64_stage_2_0_t239 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t797 = FSM_fft_64_stage_2_0_t796[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t798 = FSM_fft_64_stage_2_0_t797[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t799 = FSM_fft_64_stage_2_0_t795;
    FSM_fft_64_stage_2_0_t799[FSM_fft_64_stage_2_0_t798 * 32 +: 32] = FSM_fft_64_stage_2_0_t788 - FSM_fft_64_stage_2_0_t792;
    FSM_fft_64_stage_2_0_t800 = FSM_fft_64_stage_2_0_t273[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t801 = FSM_fft_64_stage_2_0_t273[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t802 = FSM_fft_64_stage_2_0_t799[FSM_fft_64_stage_2_0_t801 * 32 +: 32];
    FSM_fft_64_stage_2_0_t803 = FSM_fft_64_stage_2_0_t273 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t804 = FSM_fft_64_stage_2_0_t803[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t805 = FSM_fft_64_stage_2_0_t804[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t806 = FSM_fft_64_stage_2_0_t799[FSM_fft_64_stage_2_0_t805 * 32 +: 32];
    FSM_fft_64_stage_2_0_t807 = FSM_fft_64_stage_2_0_t802 + FSM_fft_64_stage_2_0_t806;
    FSM_fft_64_stage_2_0_t808 = FSM_fft_64_stage_2_0_t807[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t809 = FSM_fft_64_stage_2_0_t799;
    FSM_fft_64_stage_2_0_t809[FSM_fft_64_stage_2_0_t800 * 32 +: 32] = FSM_fft_64_stage_2_0_t808;
    FSM_fft_64_stage_2_0_t810 = FSM_fft_64_stage_2_0_t273 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t811 = FSM_fft_64_stage_2_0_t810[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t812 = FSM_fft_64_stage_2_0_t811[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t813 = FSM_fft_64_stage_2_0_t809;
    FSM_fft_64_stage_2_0_t813[FSM_fft_64_stage_2_0_t812 * 32 +: 32] = FSM_fft_64_stage_2_0_t802 - FSM_fft_64_stage_2_0_t806;
    FSM_fft_64_stage_2_0_t814 = FSM_fft_64_stage_2_0_t273 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t815 = FSM_fft_64_stage_2_0_t814[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t816 = FSM_fft_64_stage_2_0_t815[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t817 = FSM_fft_64_stage_2_0_t273 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t818 = FSM_fft_64_stage_2_0_t817[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t819 = FSM_fft_64_stage_2_0_t818[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t820 = FSM_fft_64_stage_2_0_t799[FSM_fft_64_stage_2_0_t819 * 32 +: 32];
    FSM_fft_64_stage_2_0_t821 = FSM_fft_64_stage_2_0_t273 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t822 = FSM_fft_64_stage_2_0_t821[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t823 = FSM_fft_64_stage_2_0_t822[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t824 = FSM_fft_64_stage_2_0_t799[FSM_fft_64_stage_2_0_t823 * 32 +: 32];
    FSM_fft_64_stage_2_0_t825 = FSM_fft_64_stage_2_0_t820 + FSM_fft_64_stage_2_0_t824;
    FSM_fft_64_stage_2_0_t826 = FSM_fft_64_stage_2_0_t825[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t827 = FSM_fft_64_stage_2_0_t813;
    FSM_fft_64_stage_2_0_t827[FSM_fft_64_stage_2_0_t816 * 32 +: 32] = FSM_fft_64_stage_2_0_t826;
    FSM_fft_64_stage_2_0_t828 = FSM_fft_64_stage_2_0_t273 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t829 = FSM_fft_64_stage_2_0_t828[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t830 = FSM_fft_64_stage_2_0_t829[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t831 = FSM_fft_64_stage_2_0_t827;
    FSM_fft_64_stage_2_0_t831[FSM_fft_64_stage_2_0_t830 * 32 +: 32] = FSM_fft_64_stage_2_0_t820 - FSM_fft_64_stage_2_0_t824;
    FSM_fft_64_stage_2_0_t832 = FSM_fft_64_stage_2_0_t307[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t833 = FSM_fft_64_stage_2_0_t307[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t834 = FSM_fft_64_stage_2_0_t831[FSM_fft_64_stage_2_0_t833 * 32 +: 32];
    FSM_fft_64_stage_2_0_t835 = FSM_fft_64_stage_2_0_t307 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t836 = FSM_fft_64_stage_2_0_t835[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t837 = FSM_fft_64_stage_2_0_t836[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t838 = FSM_fft_64_stage_2_0_t831[FSM_fft_64_stage_2_0_t837 * 32 +: 32];
    FSM_fft_64_stage_2_0_t839 = FSM_fft_64_stage_2_0_t834 + FSM_fft_64_stage_2_0_t838;
    FSM_fft_64_stage_2_0_t840 = FSM_fft_64_stage_2_0_t839[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t841 = FSM_fft_64_stage_2_0_t831;
    FSM_fft_64_stage_2_0_t841[FSM_fft_64_stage_2_0_t832 * 32 +: 32] = FSM_fft_64_stage_2_0_t840;
    FSM_fft_64_stage_2_0_t842 = FSM_fft_64_stage_2_0_t307 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t843 = FSM_fft_64_stage_2_0_t842[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t844 = FSM_fft_64_stage_2_0_t843[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t845 = FSM_fft_64_stage_2_0_t841;
    FSM_fft_64_stage_2_0_t845[FSM_fft_64_stage_2_0_t844 * 32 +: 32] = FSM_fft_64_stage_2_0_t834 - FSM_fft_64_stage_2_0_t838;
    FSM_fft_64_stage_2_0_t846 = FSM_fft_64_stage_2_0_t307 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t847 = FSM_fft_64_stage_2_0_t846[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t848 = FSM_fft_64_stage_2_0_t847[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t849 = FSM_fft_64_stage_2_0_t307 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t850 = FSM_fft_64_stage_2_0_t849[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t851 = FSM_fft_64_stage_2_0_t850[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t852 = FSM_fft_64_stage_2_0_t831[FSM_fft_64_stage_2_0_t851 * 32 +: 32];
    FSM_fft_64_stage_2_0_t853 = FSM_fft_64_stage_2_0_t307 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t854 = FSM_fft_64_stage_2_0_t853[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t855 = FSM_fft_64_stage_2_0_t854[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t856 = FSM_fft_64_stage_2_0_t831[FSM_fft_64_stage_2_0_t855 * 32 +: 32];
    FSM_fft_64_stage_2_0_t857 = FSM_fft_64_stage_2_0_t852 + FSM_fft_64_stage_2_0_t856;
    FSM_fft_64_stage_2_0_t858 = FSM_fft_64_stage_2_0_t857[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t859 = FSM_fft_64_stage_2_0_t845;
    FSM_fft_64_stage_2_0_t859[FSM_fft_64_stage_2_0_t848 * 32 +: 32] = FSM_fft_64_stage_2_0_t858;
    FSM_fft_64_stage_2_0_t860 = FSM_fft_64_stage_2_0_t307 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t861 = FSM_fft_64_stage_2_0_t860[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t862 = FSM_fft_64_stage_2_0_t861[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t863 = FSM_fft_64_stage_2_0_t859;
    FSM_fft_64_stage_2_0_t863[FSM_fft_64_stage_2_0_t862 * 32 +: 32] = FSM_fft_64_stage_2_0_t852 - FSM_fft_64_stage_2_0_t856;
    FSM_fft_64_stage_2_0_t864 = FSM_fft_64_stage_2_0_t341[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t865 = FSM_fft_64_stage_2_0_t341[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t866 = FSM_fft_64_stage_2_0_t863[FSM_fft_64_stage_2_0_t865 * 32 +: 32];
    FSM_fft_64_stage_2_0_t867 = FSM_fft_64_stage_2_0_t341 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t868 = FSM_fft_64_stage_2_0_t867[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t869 = FSM_fft_64_stage_2_0_t868[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t870 = FSM_fft_64_stage_2_0_t863[FSM_fft_64_stage_2_0_t869 * 32 +: 32];
    FSM_fft_64_stage_2_0_t871 = FSM_fft_64_stage_2_0_t866 + FSM_fft_64_stage_2_0_t870;
    FSM_fft_64_stage_2_0_t872 = FSM_fft_64_stage_2_0_t871[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t873 = FSM_fft_64_stage_2_0_t863;
    FSM_fft_64_stage_2_0_t873[FSM_fft_64_stage_2_0_t864 * 32 +: 32] = FSM_fft_64_stage_2_0_t872;
    FSM_fft_64_stage_2_0_t874 = FSM_fft_64_stage_2_0_t341 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t875 = FSM_fft_64_stage_2_0_t874[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t876 = FSM_fft_64_stage_2_0_t875[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t877 = FSM_fft_64_stage_2_0_t873;
    FSM_fft_64_stage_2_0_t877[FSM_fft_64_stage_2_0_t876 * 32 +: 32] = FSM_fft_64_stage_2_0_t866 - FSM_fft_64_stage_2_0_t870;
    FSM_fft_64_stage_2_0_t878 = FSM_fft_64_stage_2_0_t341 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t879 = FSM_fft_64_stage_2_0_t878[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t880 = FSM_fft_64_stage_2_0_t879[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t881 = FSM_fft_64_stage_2_0_t341 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t882 = FSM_fft_64_stage_2_0_t881[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t883 = FSM_fft_64_stage_2_0_t882[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t884 = FSM_fft_64_stage_2_0_t863[FSM_fft_64_stage_2_0_t883 * 32 +: 32];
    FSM_fft_64_stage_2_0_t885 = FSM_fft_64_stage_2_0_t341 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t886 = FSM_fft_64_stage_2_0_t885[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t887 = FSM_fft_64_stage_2_0_t886[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t888 = FSM_fft_64_stage_2_0_t863[FSM_fft_64_stage_2_0_t887 * 32 +: 32];
    FSM_fft_64_stage_2_0_t889 = FSM_fft_64_stage_2_0_t884 + FSM_fft_64_stage_2_0_t888;
    FSM_fft_64_stage_2_0_t890 = FSM_fft_64_stage_2_0_t889[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t891 = FSM_fft_64_stage_2_0_t877;
    FSM_fft_64_stage_2_0_t891[FSM_fft_64_stage_2_0_t880 * 32 +: 32] = FSM_fft_64_stage_2_0_t890;
    FSM_fft_64_stage_2_0_t892 = FSM_fft_64_stage_2_0_t341 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t893 = FSM_fft_64_stage_2_0_t892[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t894 = FSM_fft_64_stage_2_0_t893[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t895 = FSM_fft_64_stage_2_0_t891;
    FSM_fft_64_stage_2_0_t895[FSM_fft_64_stage_2_0_t894 * 32 +: 32] = FSM_fft_64_stage_2_0_t884 - FSM_fft_64_stage_2_0_t888;
    FSM_fft_64_stage_2_0_t896 = FSM_fft_64_stage_2_0_t375[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t897 = FSM_fft_64_stage_2_0_t375[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t898 = FSM_fft_64_stage_2_0_t895[FSM_fft_64_stage_2_0_t897 * 32 +: 32];
    FSM_fft_64_stage_2_0_t899 = FSM_fft_64_stage_2_0_t375 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t900 = FSM_fft_64_stage_2_0_t899[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t901 = FSM_fft_64_stage_2_0_t900[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t902 = FSM_fft_64_stage_2_0_t895[FSM_fft_64_stage_2_0_t901 * 32 +: 32];
    FSM_fft_64_stage_2_0_t903 = FSM_fft_64_stage_2_0_t898 + FSM_fft_64_stage_2_0_t902;
    FSM_fft_64_stage_2_0_t904 = FSM_fft_64_stage_2_0_t903[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t905 = FSM_fft_64_stage_2_0_t895;
    FSM_fft_64_stage_2_0_t905[FSM_fft_64_stage_2_0_t896 * 32 +: 32] = FSM_fft_64_stage_2_0_t904;
    FSM_fft_64_stage_2_0_t906 = FSM_fft_64_stage_2_0_t375 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t907 = FSM_fft_64_stage_2_0_t906[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t908 = FSM_fft_64_stage_2_0_t907[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t909 = FSM_fft_64_stage_2_0_t905;
    FSM_fft_64_stage_2_0_t909[FSM_fft_64_stage_2_0_t908 * 32 +: 32] = FSM_fft_64_stage_2_0_t898 - FSM_fft_64_stage_2_0_t902;
    FSM_fft_64_stage_2_0_t910 = FSM_fft_64_stage_2_0_t375 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t911 = FSM_fft_64_stage_2_0_t910[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t912 = FSM_fft_64_stage_2_0_t911[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t913 = FSM_fft_64_stage_2_0_t375 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t914 = FSM_fft_64_stage_2_0_t913[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t915 = FSM_fft_64_stage_2_0_t914[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t916 = FSM_fft_64_stage_2_0_t895[FSM_fft_64_stage_2_0_t915 * 32 +: 32];
    FSM_fft_64_stage_2_0_t917 = FSM_fft_64_stage_2_0_t375 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t918 = FSM_fft_64_stage_2_0_t917[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t919 = FSM_fft_64_stage_2_0_t918[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t920 = FSM_fft_64_stage_2_0_t895[FSM_fft_64_stage_2_0_t919 * 32 +: 32];
    FSM_fft_64_stage_2_0_t921 = FSM_fft_64_stage_2_0_t916 + FSM_fft_64_stage_2_0_t920;
    FSM_fft_64_stage_2_0_t922 = FSM_fft_64_stage_2_0_t921[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t923 = FSM_fft_64_stage_2_0_t909;
    FSM_fft_64_stage_2_0_t923[FSM_fft_64_stage_2_0_t912 * 32 +: 32] = FSM_fft_64_stage_2_0_t922;
    FSM_fft_64_stage_2_0_t924 = FSM_fft_64_stage_2_0_t375 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t925 = FSM_fft_64_stage_2_0_t924[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t926 = FSM_fft_64_stage_2_0_t925[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t927 = FSM_fft_64_stage_2_0_t923;
    FSM_fft_64_stage_2_0_t927[FSM_fft_64_stage_2_0_t926 * 32 +: 32] = FSM_fft_64_stage_2_0_t916 - FSM_fft_64_stage_2_0_t920;
    FSM_fft_64_stage_2_0_t928 = FSM_fft_64_stage_2_0_t409[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t929 = FSM_fft_64_stage_2_0_t409[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t930 = FSM_fft_64_stage_2_0_t927[FSM_fft_64_stage_2_0_t929 * 32 +: 32];
    FSM_fft_64_stage_2_0_t931 = FSM_fft_64_stage_2_0_t409 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t932 = FSM_fft_64_stage_2_0_t931[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t933 = FSM_fft_64_stage_2_0_t932[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t934 = FSM_fft_64_stage_2_0_t927[FSM_fft_64_stage_2_0_t933 * 32 +: 32];
    FSM_fft_64_stage_2_0_t935 = FSM_fft_64_stage_2_0_t930 + FSM_fft_64_stage_2_0_t934;
    FSM_fft_64_stage_2_0_t936 = FSM_fft_64_stage_2_0_t935[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t937 = FSM_fft_64_stage_2_0_t927;
    FSM_fft_64_stage_2_0_t937[FSM_fft_64_stage_2_0_t928 * 32 +: 32] = FSM_fft_64_stage_2_0_t936;
    FSM_fft_64_stage_2_0_t938 = FSM_fft_64_stage_2_0_t409 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t939 = FSM_fft_64_stage_2_0_t938[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t940 = FSM_fft_64_stage_2_0_t939[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t941 = FSM_fft_64_stage_2_0_t937;
    FSM_fft_64_stage_2_0_t941[FSM_fft_64_stage_2_0_t940 * 32 +: 32] = FSM_fft_64_stage_2_0_t930 - FSM_fft_64_stage_2_0_t934;
    FSM_fft_64_stage_2_0_t942 = FSM_fft_64_stage_2_0_t409 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t943 = FSM_fft_64_stage_2_0_t942[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t944 = FSM_fft_64_stage_2_0_t943[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t945 = FSM_fft_64_stage_2_0_t409 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t946 = FSM_fft_64_stage_2_0_t945[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t947 = FSM_fft_64_stage_2_0_t946[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t948 = FSM_fft_64_stage_2_0_t927[FSM_fft_64_stage_2_0_t947 * 32 +: 32];
    FSM_fft_64_stage_2_0_t949 = FSM_fft_64_stage_2_0_t409 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t950 = FSM_fft_64_stage_2_0_t949[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t951 = FSM_fft_64_stage_2_0_t950[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t952 = FSM_fft_64_stage_2_0_t927[FSM_fft_64_stage_2_0_t951 * 32 +: 32];
    FSM_fft_64_stage_2_0_t953 = FSM_fft_64_stage_2_0_t948 + FSM_fft_64_stage_2_0_t952;
    FSM_fft_64_stage_2_0_t954 = FSM_fft_64_stage_2_0_t953[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t955 = FSM_fft_64_stage_2_0_t941;
    FSM_fft_64_stage_2_0_t955[FSM_fft_64_stage_2_0_t944 * 32 +: 32] = FSM_fft_64_stage_2_0_t954;
    FSM_fft_64_stage_2_0_t956 = FSM_fft_64_stage_2_0_t409 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t957 = FSM_fft_64_stage_2_0_t956[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t958 = FSM_fft_64_stage_2_0_t957[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t959 = FSM_fft_64_stage_2_0_t955;
    FSM_fft_64_stage_2_0_t959[FSM_fft_64_stage_2_0_t958 * 32 +: 32] = FSM_fft_64_stage_2_0_t948 - FSM_fft_64_stage_2_0_t952;
    FSM_fft_64_stage_2_0_t960 = FSM_fft_64_stage_2_0_t443[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t961 = FSM_fft_64_stage_2_0_t443[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t962 = FSM_fft_64_stage_2_0_t959[FSM_fft_64_stage_2_0_t961 * 32 +: 32];
    FSM_fft_64_stage_2_0_t963 = FSM_fft_64_stage_2_0_t443 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t964 = FSM_fft_64_stage_2_0_t963[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t965 = FSM_fft_64_stage_2_0_t964[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t966 = FSM_fft_64_stage_2_0_t959[FSM_fft_64_stage_2_0_t965 * 32 +: 32];
    FSM_fft_64_stage_2_0_t967 = FSM_fft_64_stage_2_0_t962 + FSM_fft_64_stage_2_0_t966;
    FSM_fft_64_stage_2_0_t968 = FSM_fft_64_stage_2_0_t967[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t969 = FSM_fft_64_stage_2_0_t959;
    FSM_fft_64_stage_2_0_t969[FSM_fft_64_stage_2_0_t960 * 32 +: 32] = FSM_fft_64_stage_2_0_t968;
    FSM_fft_64_stage_2_0_t970 = FSM_fft_64_stage_2_0_t443 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t971 = FSM_fft_64_stage_2_0_t970[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t972 = FSM_fft_64_stage_2_0_t971[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t973 = FSM_fft_64_stage_2_0_t969;
    FSM_fft_64_stage_2_0_t973[FSM_fft_64_stage_2_0_t972 * 32 +: 32] = FSM_fft_64_stage_2_0_t962 - FSM_fft_64_stage_2_0_t966;
    FSM_fft_64_stage_2_0_t974 = FSM_fft_64_stage_2_0_t443 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t975 = FSM_fft_64_stage_2_0_t974[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t976 = FSM_fft_64_stage_2_0_t975[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t977 = FSM_fft_64_stage_2_0_t443 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t978 = FSM_fft_64_stage_2_0_t977[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t979 = FSM_fft_64_stage_2_0_t978[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t980 = FSM_fft_64_stage_2_0_t959[FSM_fft_64_stage_2_0_t979 * 32 +: 32];
    FSM_fft_64_stage_2_0_t981 = FSM_fft_64_stage_2_0_t443 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t982 = FSM_fft_64_stage_2_0_t981[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t983 = FSM_fft_64_stage_2_0_t982[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t984 = FSM_fft_64_stage_2_0_t959[FSM_fft_64_stage_2_0_t983 * 32 +: 32];
    FSM_fft_64_stage_2_0_t985 = FSM_fft_64_stage_2_0_t980 + FSM_fft_64_stage_2_0_t984;
    FSM_fft_64_stage_2_0_t986 = FSM_fft_64_stage_2_0_t985[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t987 = FSM_fft_64_stage_2_0_t973;
    FSM_fft_64_stage_2_0_t987[FSM_fft_64_stage_2_0_t976 * 32 +: 32] = FSM_fft_64_stage_2_0_t986;
    FSM_fft_64_stage_2_0_t988 = FSM_fft_64_stage_2_0_t443 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t989 = FSM_fft_64_stage_2_0_t988[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t990 = FSM_fft_64_stage_2_0_t989[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t991 = FSM_fft_64_stage_2_0_t987;
    FSM_fft_64_stage_2_0_t991[FSM_fft_64_stage_2_0_t990 * 32 +: 32] = FSM_fft_64_stage_2_0_t980 - FSM_fft_64_stage_2_0_t984;
    FSM_fft_64_stage_2_0_t992 = FSM_fft_64_stage_2_0_t477[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t993 = FSM_fft_64_stage_2_0_t477[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t994 = FSM_fft_64_stage_2_0_t991[FSM_fft_64_stage_2_0_t993 * 32 +: 32];
    FSM_fft_64_stage_2_0_t995 = FSM_fft_64_stage_2_0_t477 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t996 = FSM_fft_64_stage_2_0_t995[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t997 = FSM_fft_64_stage_2_0_t996[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t998 = FSM_fft_64_stage_2_0_t991[FSM_fft_64_stage_2_0_t997 * 32 +: 32];
    FSM_fft_64_stage_2_0_t999 = FSM_fft_64_stage_2_0_t994 + FSM_fft_64_stage_2_0_t998;
    FSM_fft_64_stage_2_0_t1000 = FSM_fft_64_stage_2_0_t999[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t1001 = FSM_fft_64_stage_2_0_t991;
    FSM_fft_64_stage_2_0_t1001[FSM_fft_64_stage_2_0_t992 * 32 +: 32] = FSM_fft_64_stage_2_0_t1000;
    FSM_fft_64_stage_2_0_t1002 = FSM_fft_64_stage_2_0_t477 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t1003 = FSM_fft_64_stage_2_0_t1002[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t1004 = FSM_fft_64_stage_2_0_t1003[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t1005 = FSM_fft_64_stage_2_0_t1001;
    FSM_fft_64_stage_2_0_t1005[FSM_fft_64_stage_2_0_t1004 * 32 +: 32] = FSM_fft_64_stage_2_0_t994 - FSM_fft_64_stage_2_0_t998;
    FSM_fft_64_stage_2_0_t1006 = FSM_fft_64_stage_2_0_t477 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t1007 = FSM_fft_64_stage_2_0_t1006[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t1008 = FSM_fft_64_stage_2_0_t1007[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t1009 = FSM_fft_64_stage_2_0_t477 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t1010 = FSM_fft_64_stage_2_0_t1009[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t1011 = FSM_fft_64_stage_2_0_t1010[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t1012 = FSM_fft_64_stage_2_0_t991[FSM_fft_64_stage_2_0_t1011 * 32 +: 32];
    FSM_fft_64_stage_2_0_t1013 = FSM_fft_64_stage_2_0_t477 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t1014 = FSM_fft_64_stage_2_0_t1013[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t1015 = FSM_fft_64_stage_2_0_t1014[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t1016 = FSM_fft_64_stage_2_0_t991[FSM_fft_64_stage_2_0_t1015 * 32 +: 32];
    FSM_fft_64_stage_2_0_t1017 = FSM_fft_64_stage_2_0_t1012 + FSM_fft_64_stage_2_0_t1016;
    FSM_fft_64_stage_2_0_t1018 = FSM_fft_64_stage_2_0_t1017[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t1019 = FSM_fft_64_stage_2_0_t1005;
    FSM_fft_64_stage_2_0_t1019[FSM_fft_64_stage_2_0_t1008 * 32 +: 32] = FSM_fft_64_stage_2_0_t1018;
    FSM_fft_64_stage_2_0_t1020 = FSM_fft_64_stage_2_0_t477 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t1021 = FSM_fft_64_stage_2_0_t1020[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t1022 = FSM_fft_64_stage_2_0_t1021[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t1023 = FSM_fft_64_stage_2_0_t1019;
    FSM_fft_64_stage_2_0_t1023[FSM_fft_64_stage_2_0_t1022 * 32 +: 32] = FSM_fft_64_stage_2_0_t1012 - FSM_fft_64_stage_2_0_t1016;
    FSM_fft_64_stage_2_0_t1024 = FSM_fft_64_stage_2_0_t511[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t1025 = FSM_fft_64_stage_2_0_t511[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t1026 = FSM_fft_64_stage_2_0_t1023[FSM_fft_64_stage_2_0_t1025 * 32 +: 32];
    FSM_fft_64_stage_2_0_t1027 = FSM_fft_64_stage_2_0_t511 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t1028 = FSM_fft_64_stage_2_0_t1027[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t1029 = FSM_fft_64_stage_2_0_t1028[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t1030 = FSM_fft_64_stage_2_0_t1023[FSM_fft_64_stage_2_0_t1029 * 32 +: 32];
    FSM_fft_64_stage_2_0_t1031 = FSM_fft_64_stage_2_0_t1026 + FSM_fft_64_stage_2_0_t1030;
    FSM_fft_64_stage_2_0_t1032 = FSM_fft_64_stage_2_0_t1031[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t1033 = FSM_fft_64_stage_2_0_t1023;
    FSM_fft_64_stage_2_0_t1033[FSM_fft_64_stage_2_0_t1024 * 32 +: 32] = FSM_fft_64_stage_2_0_t1032;
    FSM_fft_64_stage_2_0_t1034 = FSM_fft_64_stage_2_0_t511 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t1035 = FSM_fft_64_stage_2_0_t1034[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t1036 = FSM_fft_64_stage_2_0_t1035[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t1037 = FSM_fft_64_stage_2_0_t1033;
    FSM_fft_64_stage_2_0_t1037[FSM_fft_64_stage_2_0_t1036 * 32 +: 32] = FSM_fft_64_stage_2_0_t1026 - FSM_fft_64_stage_2_0_t1030;
    FSM_fft_64_stage_2_0_t1038 = FSM_fft_64_stage_2_0_t511 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t1039 = FSM_fft_64_stage_2_0_t1038[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t1040 = FSM_fft_64_stage_2_0_t1039[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t1041 = FSM_fft_64_stage_2_0_t511 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t1042 = FSM_fft_64_stage_2_0_t1041[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t1043 = FSM_fft_64_stage_2_0_t1042[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t1044 = FSM_fft_64_stage_2_0_t1023[FSM_fft_64_stage_2_0_t1043 * 32 +: 32];
    FSM_fft_64_stage_2_0_t1045 = FSM_fft_64_stage_2_0_t511 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t1046 = FSM_fft_64_stage_2_0_t1045[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t1047 = FSM_fft_64_stage_2_0_t1046[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t1048 = FSM_fft_64_stage_2_0_t1023[FSM_fft_64_stage_2_0_t1047 * 32 +: 32];
    FSM_fft_64_stage_2_0_t1049 = FSM_fft_64_stage_2_0_t1044 + FSM_fft_64_stage_2_0_t1048;
    FSM_fft_64_stage_2_0_t1050 = FSM_fft_64_stage_2_0_t1049[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t1051 = FSM_fft_64_stage_2_0_t1037;
    FSM_fft_64_stage_2_0_t1051[FSM_fft_64_stage_2_0_t1040 * 32 +: 32] = FSM_fft_64_stage_2_0_t1050;
    FSM_fft_64_stage_2_0_t1052 = FSM_fft_64_stage_2_0_t511 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t1053 = FSM_fft_64_stage_2_0_t1052[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t1054 = FSM_fft_64_stage_2_0_t1053[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t1055 = FSM_fft_64_stage_2_0_t1051;
    FSM_fft_64_stage_2_0_t1055[FSM_fft_64_stage_2_0_t1054 * 32 +: 32] = FSM_fft_64_stage_2_0_t1044 - FSM_fft_64_stage_2_0_t1048;
end

always @* begin
    FSM_fft_64_stage_2_0_t0 = 32'b0 * 32'b00000000000000000000000000000100;
    FSM_fft_64_stage_2_0_t1 = FSM_fft_64_stage_2_0_t0[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t2 = FSM_fft_64_stage_2_0_t1[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t3 = FSM_fft_64_stage_2_0_t1[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t4 = i_data_in_real[FSM_fft_64_stage_2_0_t3 * 32 +: 32];
    FSM_fft_64_stage_2_0_t5 = FSM_fft_64_stage_2_0_t1 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t6 = FSM_fft_64_stage_2_0_t5[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t7 = FSM_fft_64_stage_2_0_t6[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t8 = i_data_in_real[FSM_fft_64_stage_2_0_t7 * 32 +: 32];
    FSM_fft_64_stage_2_0_t9 = FSM_fft_64_stage_2_0_t4 + FSM_fft_64_stage_2_0_t8;
    FSM_fft_64_stage_2_0_t10 = FSM_fft_64_stage_2_0_t9[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t11 = i_data_in_real;
    FSM_fft_64_stage_2_0_t11[FSM_fft_64_stage_2_0_t2 * 32 +: 32] = FSM_fft_64_stage_2_0_t10;
    FSM_fft_64_stage_2_0_t12 = FSM_fft_64_stage_2_0_t1 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t13 = FSM_fft_64_stage_2_0_t12[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t14 = FSM_fft_64_stage_2_0_t13[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t15 = FSM_fft_64_stage_2_0_t11;
    FSM_fft_64_stage_2_0_t15[FSM_fft_64_stage_2_0_t14 * 32 +: 32] = FSM_fft_64_stage_2_0_t4 - FSM_fft_64_stage_2_0_t8;
    FSM_fft_64_stage_2_0_t16 = FSM_fft_64_stage_2_0_t1 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t17 = FSM_fft_64_stage_2_0_t16[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t18 = FSM_fft_64_stage_2_0_t17[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t19 = FSM_fft_64_stage_2_0_t1 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t20 = FSM_fft_64_stage_2_0_t19[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t21 = FSM_fft_64_stage_2_0_t20[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t22 = i_data_in_real[FSM_fft_64_stage_2_0_t21 * 32 +: 32];
    FSM_fft_64_stage_2_0_t23 = FSM_fft_64_stage_2_0_t1 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t24 = FSM_fft_64_stage_2_0_t23[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t25 = FSM_fft_64_stage_2_0_t24[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t26 = i_data_in_real[FSM_fft_64_stage_2_0_t25 * 32 +: 32];
    FSM_fft_64_stage_2_0_t27 = FSM_fft_64_stage_2_0_t22 + FSM_fft_64_stage_2_0_t26;
    FSM_fft_64_stage_2_0_t28 = FSM_fft_64_stage_2_0_t27[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t29 = FSM_fft_64_stage_2_0_t15;
    FSM_fft_64_stage_2_0_t29[FSM_fft_64_stage_2_0_t18 * 32 +: 32] = FSM_fft_64_stage_2_0_t28;
    FSM_fft_64_stage_2_0_t30 = FSM_fft_64_stage_2_0_t1 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t31 = FSM_fft_64_stage_2_0_t30[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t32 = FSM_fft_64_stage_2_0_t31[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t33 = FSM_fft_64_stage_2_0_t29;
    FSM_fft_64_stage_2_0_t33[FSM_fft_64_stage_2_0_t32 * 32 +: 32] = FSM_fft_64_stage_2_0_t22 - FSM_fft_64_stage_2_0_t26;
    FSM_fft_64_stage_2_0_t34 = 32'b00000000000000000000000000000001 * 32'b00000000000000000000000000000100;
    FSM_fft_64_stage_2_0_t35 = FSM_fft_64_stage_2_0_t34[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t36 = FSM_fft_64_stage_2_0_t35[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t37 = FSM_fft_64_stage_2_0_t35[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t38 = FSM_fft_64_stage_2_0_t33[FSM_fft_64_stage_2_0_t37 * 32 +: 32];
    FSM_fft_64_stage_2_0_t39 = FSM_fft_64_stage_2_0_t35 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t40 = FSM_fft_64_stage_2_0_t39[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t41 = FSM_fft_64_stage_2_0_t40[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t42 = FSM_fft_64_stage_2_0_t33[FSM_fft_64_stage_2_0_t41 * 32 +: 32];
    FSM_fft_64_stage_2_0_t43 = FSM_fft_64_stage_2_0_t38 + FSM_fft_64_stage_2_0_t42;
    FSM_fft_64_stage_2_0_t44 = FSM_fft_64_stage_2_0_t43[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t45 = FSM_fft_64_stage_2_0_t33;
    FSM_fft_64_stage_2_0_t45[FSM_fft_64_stage_2_0_t36 * 32 +: 32] = FSM_fft_64_stage_2_0_t44;
    FSM_fft_64_stage_2_0_t46 = FSM_fft_64_stage_2_0_t35 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t47 = FSM_fft_64_stage_2_0_t46[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t48 = FSM_fft_64_stage_2_0_t47[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t49 = FSM_fft_64_stage_2_0_t45;
    FSM_fft_64_stage_2_0_t49[FSM_fft_64_stage_2_0_t48 * 32 +: 32] = FSM_fft_64_stage_2_0_t38 - FSM_fft_64_stage_2_0_t42;
    FSM_fft_64_stage_2_0_t50 = FSM_fft_64_stage_2_0_t35 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t51 = FSM_fft_64_stage_2_0_t50[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t52 = FSM_fft_64_stage_2_0_t51[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t53 = FSM_fft_64_stage_2_0_t35 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t54 = FSM_fft_64_stage_2_0_t53[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t55 = FSM_fft_64_stage_2_0_t54[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t56 = FSM_fft_64_stage_2_0_t33[FSM_fft_64_stage_2_0_t55 * 32 +: 32];
    FSM_fft_64_stage_2_0_t57 = FSM_fft_64_stage_2_0_t35 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t58 = FSM_fft_64_stage_2_0_t57[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t59 = FSM_fft_64_stage_2_0_t58[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t60 = FSM_fft_64_stage_2_0_t33[FSM_fft_64_stage_2_0_t59 * 32 +: 32];
    FSM_fft_64_stage_2_0_t61 = FSM_fft_64_stage_2_0_t56 + FSM_fft_64_stage_2_0_t60;
    FSM_fft_64_stage_2_0_t62 = FSM_fft_64_stage_2_0_t61[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t63 = FSM_fft_64_stage_2_0_t49;
    FSM_fft_64_stage_2_0_t63[FSM_fft_64_stage_2_0_t52 * 32 +: 32] = FSM_fft_64_stage_2_0_t62;
    FSM_fft_64_stage_2_0_t64 = FSM_fft_64_stage_2_0_t35 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t65 = FSM_fft_64_stage_2_0_t64[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t66 = FSM_fft_64_stage_2_0_t65[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t67 = FSM_fft_64_stage_2_0_t63;
    FSM_fft_64_stage_2_0_t67[FSM_fft_64_stage_2_0_t66 * 32 +: 32] = FSM_fft_64_stage_2_0_t56 - FSM_fft_64_stage_2_0_t60;
    FSM_fft_64_stage_2_0_t68 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000100;
    FSM_fft_64_stage_2_0_t69 = FSM_fft_64_stage_2_0_t68[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t70 = FSM_fft_64_stage_2_0_t69[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t71 = FSM_fft_64_stage_2_0_t69[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t72 = FSM_fft_64_stage_2_0_t67[FSM_fft_64_stage_2_0_t71 * 32 +: 32];
    FSM_fft_64_stage_2_0_t73 = FSM_fft_64_stage_2_0_t69 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t74 = FSM_fft_64_stage_2_0_t73[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t75 = FSM_fft_64_stage_2_0_t74[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t76 = FSM_fft_64_stage_2_0_t67[FSM_fft_64_stage_2_0_t75 * 32 +: 32];
    FSM_fft_64_stage_2_0_t77 = FSM_fft_64_stage_2_0_t72 + FSM_fft_64_stage_2_0_t76;
    FSM_fft_64_stage_2_0_t78 = FSM_fft_64_stage_2_0_t77[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t79 = FSM_fft_64_stage_2_0_t67;
    FSM_fft_64_stage_2_0_t79[FSM_fft_64_stage_2_0_t70 * 32 +: 32] = FSM_fft_64_stage_2_0_t78;
    FSM_fft_64_stage_2_0_t80 = FSM_fft_64_stage_2_0_t69 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t81 = FSM_fft_64_stage_2_0_t80[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t82 = FSM_fft_64_stage_2_0_t81[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t83 = FSM_fft_64_stage_2_0_t79;
    FSM_fft_64_stage_2_0_t83[FSM_fft_64_stage_2_0_t82 * 32 +: 32] = FSM_fft_64_stage_2_0_t72 - FSM_fft_64_stage_2_0_t76;
    FSM_fft_64_stage_2_0_t84 = FSM_fft_64_stage_2_0_t69 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t85 = FSM_fft_64_stage_2_0_t84[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t86 = FSM_fft_64_stage_2_0_t85[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t87 = FSM_fft_64_stage_2_0_t69 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t88 = FSM_fft_64_stage_2_0_t87[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t89 = FSM_fft_64_stage_2_0_t88[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t90 = FSM_fft_64_stage_2_0_t67[FSM_fft_64_stage_2_0_t89 * 32 +: 32];
    FSM_fft_64_stage_2_0_t91 = FSM_fft_64_stage_2_0_t69 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t92 = FSM_fft_64_stage_2_0_t91[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t93 = FSM_fft_64_stage_2_0_t92[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t94 = FSM_fft_64_stage_2_0_t67[FSM_fft_64_stage_2_0_t93 * 32 +: 32];
    FSM_fft_64_stage_2_0_t95 = FSM_fft_64_stage_2_0_t90 + FSM_fft_64_stage_2_0_t94;
    FSM_fft_64_stage_2_0_t96 = FSM_fft_64_stage_2_0_t95[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t97 = FSM_fft_64_stage_2_0_t83;
    FSM_fft_64_stage_2_0_t97[FSM_fft_64_stage_2_0_t86 * 32 +: 32] = FSM_fft_64_stage_2_0_t96;
    FSM_fft_64_stage_2_0_t98 = FSM_fft_64_stage_2_0_t69 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t99 = FSM_fft_64_stage_2_0_t98[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t100 = FSM_fft_64_stage_2_0_t99[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t101 = FSM_fft_64_stage_2_0_t97;
    FSM_fft_64_stage_2_0_t101[FSM_fft_64_stage_2_0_t100 * 32 +: 32] = FSM_fft_64_stage_2_0_t90 - FSM_fft_64_stage_2_0_t94;
    FSM_fft_64_stage_2_0_t102 = 32'b00000000000000000000000000000011 * 32'b00000000000000000000000000000100;
    FSM_fft_64_stage_2_0_t103 = FSM_fft_64_stage_2_0_t102[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t104 = FSM_fft_64_stage_2_0_t103[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t105 = FSM_fft_64_stage_2_0_t103[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t106 = FSM_fft_64_stage_2_0_t101[FSM_fft_64_stage_2_0_t105 * 32 +: 32];
    FSM_fft_64_stage_2_0_t107 = FSM_fft_64_stage_2_0_t103 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t108 = FSM_fft_64_stage_2_0_t107[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t109 = FSM_fft_64_stage_2_0_t108[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t110 = FSM_fft_64_stage_2_0_t101[FSM_fft_64_stage_2_0_t109 * 32 +: 32];
    FSM_fft_64_stage_2_0_t111 = FSM_fft_64_stage_2_0_t106 + FSM_fft_64_stage_2_0_t110;
    FSM_fft_64_stage_2_0_t112 = FSM_fft_64_stage_2_0_t111[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t113 = FSM_fft_64_stage_2_0_t101;
    FSM_fft_64_stage_2_0_t113[FSM_fft_64_stage_2_0_t104 * 32 +: 32] = FSM_fft_64_stage_2_0_t112;
    FSM_fft_64_stage_2_0_t114 = FSM_fft_64_stage_2_0_t103 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t115 = FSM_fft_64_stage_2_0_t114[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t116 = FSM_fft_64_stage_2_0_t115[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t117 = FSM_fft_64_stage_2_0_t113;
    FSM_fft_64_stage_2_0_t117[FSM_fft_64_stage_2_0_t116 * 32 +: 32] = FSM_fft_64_stage_2_0_t106 - FSM_fft_64_stage_2_0_t110;
    FSM_fft_64_stage_2_0_t118 = FSM_fft_64_stage_2_0_t103 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t119 = FSM_fft_64_stage_2_0_t118[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t120 = FSM_fft_64_stage_2_0_t119[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t121 = FSM_fft_64_stage_2_0_t103 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t122 = FSM_fft_64_stage_2_0_t121[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t123 = FSM_fft_64_stage_2_0_t122[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t124 = FSM_fft_64_stage_2_0_t101[FSM_fft_64_stage_2_0_t123 * 32 +: 32];
    FSM_fft_64_stage_2_0_t125 = FSM_fft_64_stage_2_0_t103 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t126 = FSM_fft_64_stage_2_0_t125[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t127 = FSM_fft_64_stage_2_0_t126[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t128 = FSM_fft_64_stage_2_0_t101[FSM_fft_64_stage_2_0_t127 * 32 +: 32];
    FSM_fft_64_stage_2_0_t129 = FSM_fft_64_stage_2_0_t124 + FSM_fft_64_stage_2_0_t128;
    FSM_fft_64_stage_2_0_t130 = FSM_fft_64_stage_2_0_t129[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t131 = FSM_fft_64_stage_2_0_t117;
    FSM_fft_64_stage_2_0_t131[FSM_fft_64_stage_2_0_t120 * 32 +: 32] = FSM_fft_64_stage_2_0_t130;
    FSM_fft_64_stage_2_0_t132 = FSM_fft_64_stage_2_0_t103 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t133 = FSM_fft_64_stage_2_0_t132[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t134 = FSM_fft_64_stage_2_0_t133[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t135 = FSM_fft_64_stage_2_0_t131;
    FSM_fft_64_stage_2_0_t135[FSM_fft_64_stage_2_0_t134 * 32 +: 32] = FSM_fft_64_stage_2_0_t124 - FSM_fft_64_stage_2_0_t128;
    FSM_fft_64_stage_2_0_t136 = 32'b00000000000000000000000000000100 * 32'b00000000000000000000000000000100;
    FSM_fft_64_stage_2_0_t137 = FSM_fft_64_stage_2_0_t136[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t138 = FSM_fft_64_stage_2_0_t137[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t139 = FSM_fft_64_stage_2_0_t137[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t140 = FSM_fft_64_stage_2_0_t135[FSM_fft_64_stage_2_0_t139 * 32 +: 32];
    FSM_fft_64_stage_2_0_t141 = FSM_fft_64_stage_2_0_t137 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t142 = FSM_fft_64_stage_2_0_t141[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t143 = FSM_fft_64_stage_2_0_t142[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t144 = FSM_fft_64_stage_2_0_t135[FSM_fft_64_stage_2_0_t143 * 32 +: 32];
    FSM_fft_64_stage_2_0_t145 = FSM_fft_64_stage_2_0_t140 + FSM_fft_64_stage_2_0_t144;
    FSM_fft_64_stage_2_0_t146 = FSM_fft_64_stage_2_0_t145[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t147 = FSM_fft_64_stage_2_0_t135;
    FSM_fft_64_stage_2_0_t147[FSM_fft_64_stage_2_0_t138 * 32 +: 32] = FSM_fft_64_stage_2_0_t146;
    FSM_fft_64_stage_2_0_t148 = FSM_fft_64_stage_2_0_t137 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t149 = FSM_fft_64_stage_2_0_t148[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t150 = FSM_fft_64_stage_2_0_t149[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t151 = FSM_fft_64_stage_2_0_t147;
    FSM_fft_64_stage_2_0_t151[FSM_fft_64_stage_2_0_t150 * 32 +: 32] = FSM_fft_64_stage_2_0_t140 - FSM_fft_64_stage_2_0_t144;
    FSM_fft_64_stage_2_0_t152 = FSM_fft_64_stage_2_0_t137 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t153 = FSM_fft_64_stage_2_0_t152[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t154 = FSM_fft_64_stage_2_0_t153[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t155 = FSM_fft_64_stage_2_0_t137 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t156 = FSM_fft_64_stage_2_0_t155[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t157 = FSM_fft_64_stage_2_0_t156[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t158 = FSM_fft_64_stage_2_0_t135[FSM_fft_64_stage_2_0_t157 * 32 +: 32];
    FSM_fft_64_stage_2_0_t159 = FSM_fft_64_stage_2_0_t137 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t160 = FSM_fft_64_stage_2_0_t159[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t161 = FSM_fft_64_stage_2_0_t160[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t162 = FSM_fft_64_stage_2_0_t135[FSM_fft_64_stage_2_0_t161 * 32 +: 32];
    FSM_fft_64_stage_2_0_t163 = FSM_fft_64_stage_2_0_t158 + FSM_fft_64_stage_2_0_t162;
    FSM_fft_64_stage_2_0_t164 = FSM_fft_64_stage_2_0_t163[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t165 = FSM_fft_64_stage_2_0_t151;
    FSM_fft_64_stage_2_0_t165[FSM_fft_64_stage_2_0_t154 * 32 +: 32] = FSM_fft_64_stage_2_0_t164;
    FSM_fft_64_stage_2_0_t166 = FSM_fft_64_stage_2_0_t137 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t167 = FSM_fft_64_stage_2_0_t166[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t168 = FSM_fft_64_stage_2_0_t167[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t169 = FSM_fft_64_stage_2_0_t165;
    FSM_fft_64_stage_2_0_t169[FSM_fft_64_stage_2_0_t168 * 32 +: 32] = FSM_fft_64_stage_2_0_t158 - FSM_fft_64_stage_2_0_t162;
    FSM_fft_64_stage_2_0_t170 = 32'b00000000000000000000000000000101 * 32'b00000000000000000000000000000100;
    FSM_fft_64_stage_2_0_t171 = FSM_fft_64_stage_2_0_t170[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t172 = FSM_fft_64_stage_2_0_t171[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t173 = FSM_fft_64_stage_2_0_t171[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t174 = FSM_fft_64_stage_2_0_t169[FSM_fft_64_stage_2_0_t173 * 32 +: 32];
    FSM_fft_64_stage_2_0_t175 = FSM_fft_64_stage_2_0_t171 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t176 = FSM_fft_64_stage_2_0_t175[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t177 = FSM_fft_64_stage_2_0_t176[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t178 = FSM_fft_64_stage_2_0_t169[FSM_fft_64_stage_2_0_t177 * 32 +: 32];
    FSM_fft_64_stage_2_0_t179 = FSM_fft_64_stage_2_0_t174 + FSM_fft_64_stage_2_0_t178;
    FSM_fft_64_stage_2_0_t180 = FSM_fft_64_stage_2_0_t179[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t181 = FSM_fft_64_stage_2_0_t169;
    FSM_fft_64_stage_2_0_t181[FSM_fft_64_stage_2_0_t172 * 32 +: 32] = FSM_fft_64_stage_2_0_t180;
    FSM_fft_64_stage_2_0_t182 = FSM_fft_64_stage_2_0_t171 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t183 = FSM_fft_64_stage_2_0_t182[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t184 = FSM_fft_64_stage_2_0_t183[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t185 = FSM_fft_64_stage_2_0_t181;
    FSM_fft_64_stage_2_0_t185[FSM_fft_64_stage_2_0_t184 * 32 +: 32] = FSM_fft_64_stage_2_0_t174 - FSM_fft_64_stage_2_0_t178;
    FSM_fft_64_stage_2_0_t186 = FSM_fft_64_stage_2_0_t171 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t187 = FSM_fft_64_stage_2_0_t186[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t188 = FSM_fft_64_stage_2_0_t187[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t189 = FSM_fft_64_stage_2_0_t171 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t190 = FSM_fft_64_stage_2_0_t189[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t191 = FSM_fft_64_stage_2_0_t190[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t192 = FSM_fft_64_stage_2_0_t169[FSM_fft_64_stage_2_0_t191 * 32 +: 32];
    FSM_fft_64_stage_2_0_t193 = FSM_fft_64_stage_2_0_t171 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t194 = FSM_fft_64_stage_2_0_t193[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t195 = FSM_fft_64_stage_2_0_t194[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t196 = FSM_fft_64_stage_2_0_t169[FSM_fft_64_stage_2_0_t195 * 32 +: 32];
    FSM_fft_64_stage_2_0_t197 = FSM_fft_64_stage_2_0_t192 + FSM_fft_64_stage_2_0_t196;
    FSM_fft_64_stage_2_0_t198 = FSM_fft_64_stage_2_0_t197[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t199 = FSM_fft_64_stage_2_0_t185;
    FSM_fft_64_stage_2_0_t199[FSM_fft_64_stage_2_0_t188 * 32 +: 32] = FSM_fft_64_stage_2_0_t198;
    FSM_fft_64_stage_2_0_t200 = FSM_fft_64_stage_2_0_t171 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t201 = FSM_fft_64_stage_2_0_t200[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t202 = FSM_fft_64_stage_2_0_t201[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t203 = FSM_fft_64_stage_2_0_t199;
    FSM_fft_64_stage_2_0_t203[FSM_fft_64_stage_2_0_t202 * 32 +: 32] = FSM_fft_64_stage_2_0_t192 - FSM_fft_64_stage_2_0_t196;
    FSM_fft_64_stage_2_0_t204 = 32'b00000000000000000000000000000110 * 32'b00000000000000000000000000000100;
    FSM_fft_64_stage_2_0_t205 = FSM_fft_64_stage_2_0_t204[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t206 = FSM_fft_64_stage_2_0_t205[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t207 = FSM_fft_64_stage_2_0_t205[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t208 = FSM_fft_64_stage_2_0_t203[FSM_fft_64_stage_2_0_t207 * 32 +: 32];
    FSM_fft_64_stage_2_0_t209 = FSM_fft_64_stage_2_0_t205 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t210 = FSM_fft_64_stage_2_0_t209[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t211 = FSM_fft_64_stage_2_0_t210[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t212 = FSM_fft_64_stage_2_0_t203[FSM_fft_64_stage_2_0_t211 * 32 +: 32];
    FSM_fft_64_stage_2_0_t213 = FSM_fft_64_stage_2_0_t208 + FSM_fft_64_stage_2_0_t212;
    FSM_fft_64_stage_2_0_t214 = FSM_fft_64_stage_2_0_t213[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t215 = FSM_fft_64_stage_2_0_t203;
    FSM_fft_64_stage_2_0_t215[FSM_fft_64_stage_2_0_t206 * 32 +: 32] = FSM_fft_64_stage_2_0_t214;
    FSM_fft_64_stage_2_0_t216 = FSM_fft_64_stage_2_0_t205 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t217 = FSM_fft_64_stage_2_0_t216[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t218 = FSM_fft_64_stage_2_0_t217[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t219 = FSM_fft_64_stage_2_0_t215;
    FSM_fft_64_stage_2_0_t219[FSM_fft_64_stage_2_0_t218 * 32 +: 32] = FSM_fft_64_stage_2_0_t208 - FSM_fft_64_stage_2_0_t212;
    FSM_fft_64_stage_2_0_t220 = FSM_fft_64_stage_2_0_t205 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t221 = FSM_fft_64_stage_2_0_t220[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t222 = FSM_fft_64_stage_2_0_t221[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t223 = FSM_fft_64_stage_2_0_t205 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t224 = FSM_fft_64_stage_2_0_t223[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t225 = FSM_fft_64_stage_2_0_t224[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t226 = FSM_fft_64_stage_2_0_t203[FSM_fft_64_stage_2_0_t225 * 32 +: 32];
    FSM_fft_64_stage_2_0_t227 = FSM_fft_64_stage_2_0_t205 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t228 = FSM_fft_64_stage_2_0_t227[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t229 = FSM_fft_64_stage_2_0_t228[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t230 = FSM_fft_64_stage_2_0_t203[FSM_fft_64_stage_2_0_t229 * 32 +: 32];
    FSM_fft_64_stage_2_0_t231 = FSM_fft_64_stage_2_0_t226 + FSM_fft_64_stage_2_0_t230;
    FSM_fft_64_stage_2_0_t232 = FSM_fft_64_stage_2_0_t231[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t233 = FSM_fft_64_stage_2_0_t219;
    FSM_fft_64_stage_2_0_t233[FSM_fft_64_stage_2_0_t222 * 32 +: 32] = FSM_fft_64_stage_2_0_t232;
    FSM_fft_64_stage_2_0_t234 = FSM_fft_64_stage_2_0_t205 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t235 = FSM_fft_64_stage_2_0_t234[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t236 = FSM_fft_64_stage_2_0_t235[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t237 = FSM_fft_64_stage_2_0_t233;
    FSM_fft_64_stage_2_0_t237[FSM_fft_64_stage_2_0_t236 * 32 +: 32] = FSM_fft_64_stage_2_0_t226 - FSM_fft_64_stage_2_0_t230;
    FSM_fft_64_stage_2_0_t238 = 32'b00000000000000000000000000000111 * 32'b00000000000000000000000000000100;
    FSM_fft_64_stage_2_0_t239 = FSM_fft_64_stage_2_0_t238[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t240 = FSM_fft_64_stage_2_0_t239[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t241 = FSM_fft_64_stage_2_0_t239[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t242 = FSM_fft_64_stage_2_0_t237[FSM_fft_64_stage_2_0_t241 * 32 +: 32];
    FSM_fft_64_stage_2_0_t243 = FSM_fft_64_stage_2_0_t239 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t244 = FSM_fft_64_stage_2_0_t243[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t245 = FSM_fft_64_stage_2_0_t244[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t246 = FSM_fft_64_stage_2_0_t237[FSM_fft_64_stage_2_0_t245 * 32 +: 32];
    FSM_fft_64_stage_2_0_t247 = FSM_fft_64_stage_2_0_t242 + FSM_fft_64_stage_2_0_t246;
    FSM_fft_64_stage_2_0_t248 = FSM_fft_64_stage_2_0_t247[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t249 = FSM_fft_64_stage_2_0_t237;
    FSM_fft_64_stage_2_0_t249[FSM_fft_64_stage_2_0_t240 * 32 +: 32] = FSM_fft_64_stage_2_0_t248;
    FSM_fft_64_stage_2_0_t250 = FSM_fft_64_stage_2_0_t239 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t251 = FSM_fft_64_stage_2_0_t250[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t252 = FSM_fft_64_stage_2_0_t251[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t253 = FSM_fft_64_stage_2_0_t249;
    FSM_fft_64_stage_2_0_t253[FSM_fft_64_stage_2_0_t252 * 32 +: 32] = FSM_fft_64_stage_2_0_t242 - FSM_fft_64_stage_2_0_t246;
    FSM_fft_64_stage_2_0_t254 = FSM_fft_64_stage_2_0_t239 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t255 = FSM_fft_64_stage_2_0_t254[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t256 = FSM_fft_64_stage_2_0_t255[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t257 = FSM_fft_64_stage_2_0_t239 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t258 = FSM_fft_64_stage_2_0_t257[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t259 = FSM_fft_64_stage_2_0_t258[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t260 = FSM_fft_64_stage_2_0_t237[FSM_fft_64_stage_2_0_t259 * 32 +: 32];
    FSM_fft_64_stage_2_0_t261 = FSM_fft_64_stage_2_0_t239 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t262 = FSM_fft_64_stage_2_0_t261[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t263 = FSM_fft_64_stage_2_0_t262[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t264 = FSM_fft_64_stage_2_0_t237[FSM_fft_64_stage_2_0_t263 * 32 +: 32];
    FSM_fft_64_stage_2_0_t265 = FSM_fft_64_stage_2_0_t260 + FSM_fft_64_stage_2_0_t264;
    FSM_fft_64_stage_2_0_t266 = FSM_fft_64_stage_2_0_t265[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t267 = FSM_fft_64_stage_2_0_t253;
    FSM_fft_64_stage_2_0_t267[FSM_fft_64_stage_2_0_t256 * 32 +: 32] = FSM_fft_64_stage_2_0_t266;
    FSM_fft_64_stage_2_0_t268 = FSM_fft_64_stage_2_0_t239 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t269 = FSM_fft_64_stage_2_0_t268[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t270 = FSM_fft_64_stage_2_0_t269[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t271 = FSM_fft_64_stage_2_0_t267;
    FSM_fft_64_stage_2_0_t271[FSM_fft_64_stage_2_0_t270 * 32 +: 32] = FSM_fft_64_stage_2_0_t260 - FSM_fft_64_stage_2_0_t264;
    FSM_fft_64_stage_2_0_t272 = 32'b00000000000000000000000000001000 * 32'b00000000000000000000000000000100;
    FSM_fft_64_stage_2_0_t273 = FSM_fft_64_stage_2_0_t272[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t274 = FSM_fft_64_stage_2_0_t273[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t275 = FSM_fft_64_stage_2_0_t273[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t276 = FSM_fft_64_stage_2_0_t271[FSM_fft_64_stage_2_0_t275 * 32 +: 32];
    FSM_fft_64_stage_2_0_t277 = FSM_fft_64_stage_2_0_t273 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t278 = FSM_fft_64_stage_2_0_t277[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t279 = FSM_fft_64_stage_2_0_t278[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t280 = FSM_fft_64_stage_2_0_t271[FSM_fft_64_stage_2_0_t279 * 32 +: 32];
    FSM_fft_64_stage_2_0_t281 = FSM_fft_64_stage_2_0_t276 + FSM_fft_64_stage_2_0_t280;
    FSM_fft_64_stage_2_0_t282 = FSM_fft_64_stage_2_0_t281[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t283 = FSM_fft_64_stage_2_0_t271;
    FSM_fft_64_stage_2_0_t283[FSM_fft_64_stage_2_0_t274 * 32 +: 32] = FSM_fft_64_stage_2_0_t282;
    FSM_fft_64_stage_2_0_t284 = FSM_fft_64_stage_2_0_t273 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t285 = FSM_fft_64_stage_2_0_t284[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t286 = FSM_fft_64_stage_2_0_t285[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t287 = FSM_fft_64_stage_2_0_t283;
    FSM_fft_64_stage_2_0_t287[FSM_fft_64_stage_2_0_t286 * 32 +: 32] = FSM_fft_64_stage_2_0_t276 - FSM_fft_64_stage_2_0_t280;
    FSM_fft_64_stage_2_0_t288 = FSM_fft_64_stage_2_0_t273 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t289 = FSM_fft_64_stage_2_0_t288[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t290 = FSM_fft_64_stage_2_0_t289[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t291 = FSM_fft_64_stage_2_0_t273 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t292 = FSM_fft_64_stage_2_0_t291[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t293 = FSM_fft_64_stage_2_0_t292[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t294 = FSM_fft_64_stage_2_0_t271[FSM_fft_64_stage_2_0_t293 * 32 +: 32];
    FSM_fft_64_stage_2_0_t295 = FSM_fft_64_stage_2_0_t273 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t296 = FSM_fft_64_stage_2_0_t295[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t297 = FSM_fft_64_stage_2_0_t296[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t298 = FSM_fft_64_stage_2_0_t271[FSM_fft_64_stage_2_0_t297 * 32 +: 32];
    FSM_fft_64_stage_2_0_t299 = FSM_fft_64_stage_2_0_t294 + FSM_fft_64_stage_2_0_t298;
    FSM_fft_64_stage_2_0_t300 = FSM_fft_64_stage_2_0_t299[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t301 = FSM_fft_64_stage_2_0_t287;
    FSM_fft_64_stage_2_0_t301[FSM_fft_64_stage_2_0_t290 * 32 +: 32] = FSM_fft_64_stage_2_0_t300;
    FSM_fft_64_stage_2_0_t302 = FSM_fft_64_stage_2_0_t273 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t303 = FSM_fft_64_stage_2_0_t302[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t304 = FSM_fft_64_stage_2_0_t303[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t305 = FSM_fft_64_stage_2_0_t301;
    FSM_fft_64_stage_2_0_t305[FSM_fft_64_stage_2_0_t304 * 32 +: 32] = FSM_fft_64_stage_2_0_t294 - FSM_fft_64_stage_2_0_t298;
    FSM_fft_64_stage_2_0_t306 = 32'b00000000000000000000000000001001 * 32'b00000000000000000000000000000100;
    FSM_fft_64_stage_2_0_t307 = FSM_fft_64_stage_2_0_t306[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t308 = FSM_fft_64_stage_2_0_t307[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t309 = FSM_fft_64_stage_2_0_t307[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t310 = FSM_fft_64_stage_2_0_t305[FSM_fft_64_stage_2_0_t309 * 32 +: 32];
    FSM_fft_64_stage_2_0_t311 = FSM_fft_64_stage_2_0_t307 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t312 = FSM_fft_64_stage_2_0_t311[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t313 = FSM_fft_64_stage_2_0_t312[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t314 = FSM_fft_64_stage_2_0_t305[FSM_fft_64_stage_2_0_t313 * 32 +: 32];
    FSM_fft_64_stage_2_0_t315 = FSM_fft_64_stage_2_0_t310 + FSM_fft_64_stage_2_0_t314;
    FSM_fft_64_stage_2_0_t316 = FSM_fft_64_stage_2_0_t315[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t317 = FSM_fft_64_stage_2_0_t305;
    FSM_fft_64_stage_2_0_t317[FSM_fft_64_stage_2_0_t308 * 32 +: 32] = FSM_fft_64_stage_2_0_t316;
    FSM_fft_64_stage_2_0_t318 = FSM_fft_64_stage_2_0_t307 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t319 = FSM_fft_64_stage_2_0_t318[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t320 = FSM_fft_64_stage_2_0_t319[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t321 = FSM_fft_64_stage_2_0_t317;
    FSM_fft_64_stage_2_0_t321[FSM_fft_64_stage_2_0_t320 * 32 +: 32] = FSM_fft_64_stage_2_0_t310 - FSM_fft_64_stage_2_0_t314;
    FSM_fft_64_stage_2_0_t322 = FSM_fft_64_stage_2_0_t307 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t323 = FSM_fft_64_stage_2_0_t322[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t324 = FSM_fft_64_stage_2_0_t323[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t325 = FSM_fft_64_stage_2_0_t307 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t326 = FSM_fft_64_stage_2_0_t325[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t327 = FSM_fft_64_stage_2_0_t326[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t328 = FSM_fft_64_stage_2_0_t305[FSM_fft_64_stage_2_0_t327 * 32 +: 32];
    FSM_fft_64_stage_2_0_t329 = FSM_fft_64_stage_2_0_t307 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t330 = FSM_fft_64_stage_2_0_t329[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t331 = FSM_fft_64_stage_2_0_t330[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t332 = FSM_fft_64_stage_2_0_t305[FSM_fft_64_stage_2_0_t331 * 32 +: 32];
    FSM_fft_64_stage_2_0_t333 = FSM_fft_64_stage_2_0_t328 + FSM_fft_64_stage_2_0_t332;
    FSM_fft_64_stage_2_0_t334 = FSM_fft_64_stage_2_0_t333[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t335 = FSM_fft_64_stage_2_0_t321;
    FSM_fft_64_stage_2_0_t335[FSM_fft_64_stage_2_0_t324 * 32 +: 32] = FSM_fft_64_stage_2_0_t334;
    FSM_fft_64_stage_2_0_t336 = FSM_fft_64_stage_2_0_t307 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t337 = FSM_fft_64_stage_2_0_t336[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t338 = FSM_fft_64_stage_2_0_t337[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t339 = FSM_fft_64_stage_2_0_t335;
    FSM_fft_64_stage_2_0_t339[FSM_fft_64_stage_2_0_t338 * 32 +: 32] = FSM_fft_64_stage_2_0_t328 - FSM_fft_64_stage_2_0_t332;
    FSM_fft_64_stage_2_0_t340 = 32'b00000000000000000000000000001010 * 32'b00000000000000000000000000000100;
    FSM_fft_64_stage_2_0_t341 = FSM_fft_64_stage_2_0_t340[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t342 = FSM_fft_64_stage_2_0_t341[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t343 = FSM_fft_64_stage_2_0_t341[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t344 = FSM_fft_64_stage_2_0_t339[FSM_fft_64_stage_2_0_t343 * 32 +: 32];
    FSM_fft_64_stage_2_0_t345 = FSM_fft_64_stage_2_0_t341 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t346 = FSM_fft_64_stage_2_0_t345[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t347 = FSM_fft_64_stage_2_0_t346[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t348 = FSM_fft_64_stage_2_0_t339[FSM_fft_64_stage_2_0_t347 * 32 +: 32];
    FSM_fft_64_stage_2_0_t349 = FSM_fft_64_stage_2_0_t344 + FSM_fft_64_stage_2_0_t348;
    FSM_fft_64_stage_2_0_t350 = FSM_fft_64_stage_2_0_t349[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t351 = FSM_fft_64_stage_2_0_t339;
    FSM_fft_64_stage_2_0_t351[FSM_fft_64_stage_2_0_t342 * 32 +: 32] = FSM_fft_64_stage_2_0_t350;
    FSM_fft_64_stage_2_0_t352 = FSM_fft_64_stage_2_0_t341 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t353 = FSM_fft_64_stage_2_0_t352[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t354 = FSM_fft_64_stage_2_0_t353[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t355 = FSM_fft_64_stage_2_0_t351;
    FSM_fft_64_stage_2_0_t355[FSM_fft_64_stage_2_0_t354 * 32 +: 32] = FSM_fft_64_stage_2_0_t344 - FSM_fft_64_stage_2_0_t348;
    FSM_fft_64_stage_2_0_t356 = FSM_fft_64_stage_2_0_t341 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t357 = FSM_fft_64_stage_2_0_t356[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t358 = FSM_fft_64_stage_2_0_t357[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t359 = FSM_fft_64_stage_2_0_t341 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t360 = FSM_fft_64_stage_2_0_t359[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t361 = FSM_fft_64_stage_2_0_t360[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t362 = FSM_fft_64_stage_2_0_t339[FSM_fft_64_stage_2_0_t361 * 32 +: 32];
    FSM_fft_64_stage_2_0_t363 = FSM_fft_64_stage_2_0_t341 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t364 = FSM_fft_64_stage_2_0_t363[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t365 = FSM_fft_64_stage_2_0_t364[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t366 = FSM_fft_64_stage_2_0_t339[FSM_fft_64_stage_2_0_t365 * 32 +: 32];
    FSM_fft_64_stage_2_0_t367 = FSM_fft_64_stage_2_0_t362 + FSM_fft_64_stage_2_0_t366;
    FSM_fft_64_stage_2_0_t368 = FSM_fft_64_stage_2_0_t367[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t369 = FSM_fft_64_stage_2_0_t355;
    FSM_fft_64_stage_2_0_t369[FSM_fft_64_stage_2_0_t358 * 32 +: 32] = FSM_fft_64_stage_2_0_t368;
    FSM_fft_64_stage_2_0_t370 = FSM_fft_64_stage_2_0_t341 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t371 = FSM_fft_64_stage_2_0_t370[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t372 = FSM_fft_64_stage_2_0_t371[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t373 = FSM_fft_64_stage_2_0_t369;
    FSM_fft_64_stage_2_0_t373[FSM_fft_64_stage_2_0_t372 * 32 +: 32] = FSM_fft_64_stage_2_0_t362 - FSM_fft_64_stage_2_0_t366;
    FSM_fft_64_stage_2_0_t374 = 32'b00000000000000000000000000001011 * 32'b00000000000000000000000000000100;
    FSM_fft_64_stage_2_0_t375 = FSM_fft_64_stage_2_0_t374[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t376 = FSM_fft_64_stage_2_0_t375[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t377 = FSM_fft_64_stage_2_0_t375[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t378 = FSM_fft_64_stage_2_0_t373[FSM_fft_64_stage_2_0_t377 * 32 +: 32];
    FSM_fft_64_stage_2_0_t379 = FSM_fft_64_stage_2_0_t375 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t380 = FSM_fft_64_stage_2_0_t379[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t381 = FSM_fft_64_stage_2_0_t380[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t382 = FSM_fft_64_stage_2_0_t373[FSM_fft_64_stage_2_0_t381 * 32 +: 32];
    FSM_fft_64_stage_2_0_t383 = FSM_fft_64_stage_2_0_t378 + FSM_fft_64_stage_2_0_t382;
    FSM_fft_64_stage_2_0_t384 = FSM_fft_64_stage_2_0_t383[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t385 = FSM_fft_64_stage_2_0_t373;
    FSM_fft_64_stage_2_0_t385[FSM_fft_64_stage_2_0_t376 * 32 +: 32] = FSM_fft_64_stage_2_0_t384;
    FSM_fft_64_stage_2_0_t386 = FSM_fft_64_stage_2_0_t375 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t387 = FSM_fft_64_stage_2_0_t386[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t388 = FSM_fft_64_stage_2_0_t387[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t389 = FSM_fft_64_stage_2_0_t385;
    FSM_fft_64_stage_2_0_t389[FSM_fft_64_stage_2_0_t388 * 32 +: 32] = FSM_fft_64_stage_2_0_t378 - FSM_fft_64_stage_2_0_t382;
    FSM_fft_64_stage_2_0_t390 = FSM_fft_64_stage_2_0_t375 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t391 = FSM_fft_64_stage_2_0_t390[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t392 = FSM_fft_64_stage_2_0_t391[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t393 = FSM_fft_64_stage_2_0_t375 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t394 = FSM_fft_64_stage_2_0_t393[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t395 = FSM_fft_64_stage_2_0_t394[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t396 = FSM_fft_64_stage_2_0_t373[FSM_fft_64_stage_2_0_t395 * 32 +: 32];
    FSM_fft_64_stage_2_0_t397 = FSM_fft_64_stage_2_0_t375 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t398 = FSM_fft_64_stage_2_0_t397[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t399 = FSM_fft_64_stage_2_0_t398[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t400 = FSM_fft_64_stage_2_0_t373[FSM_fft_64_stage_2_0_t399 * 32 +: 32];
    FSM_fft_64_stage_2_0_t401 = FSM_fft_64_stage_2_0_t396 + FSM_fft_64_stage_2_0_t400;
    FSM_fft_64_stage_2_0_t402 = FSM_fft_64_stage_2_0_t401[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t403 = FSM_fft_64_stage_2_0_t389;
    FSM_fft_64_stage_2_0_t403[FSM_fft_64_stage_2_0_t392 * 32 +: 32] = FSM_fft_64_stage_2_0_t402;
    FSM_fft_64_stage_2_0_t404 = FSM_fft_64_stage_2_0_t375 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t405 = FSM_fft_64_stage_2_0_t404[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t406 = FSM_fft_64_stage_2_0_t405[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t407 = FSM_fft_64_stage_2_0_t403;
    FSM_fft_64_stage_2_0_t407[FSM_fft_64_stage_2_0_t406 * 32 +: 32] = FSM_fft_64_stage_2_0_t396 - FSM_fft_64_stage_2_0_t400;
    FSM_fft_64_stage_2_0_t408 = 32'b00000000000000000000000000001100 * 32'b00000000000000000000000000000100;
    FSM_fft_64_stage_2_0_t409 = FSM_fft_64_stage_2_0_t408[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t410 = FSM_fft_64_stage_2_0_t409[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t411 = FSM_fft_64_stage_2_0_t409[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t412 = FSM_fft_64_stage_2_0_t407[FSM_fft_64_stage_2_0_t411 * 32 +: 32];
    FSM_fft_64_stage_2_0_t413 = FSM_fft_64_stage_2_0_t409 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t414 = FSM_fft_64_stage_2_0_t413[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t415 = FSM_fft_64_stage_2_0_t414[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t416 = FSM_fft_64_stage_2_0_t407[FSM_fft_64_stage_2_0_t415 * 32 +: 32];
    FSM_fft_64_stage_2_0_t417 = FSM_fft_64_stage_2_0_t412 + FSM_fft_64_stage_2_0_t416;
    FSM_fft_64_stage_2_0_t418 = FSM_fft_64_stage_2_0_t417[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t419 = FSM_fft_64_stage_2_0_t407;
    FSM_fft_64_stage_2_0_t419[FSM_fft_64_stage_2_0_t410 * 32 +: 32] = FSM_fft_64_stage_2_0_t418;
    FSM_fft_64_stage_2_0_t420 = FSM_fft_64_stage_2_0_t409 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t421 = FSM_fft_64_stage_2_0_t420[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t422 = FSM_fft_64_stage_2_0_t421[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t423 = FSM_fft_64_stage_2_0_t419;
    FSM_fft_64_stage_2_0_t423[FSM_fft_64_stage_2_0_t422 * 32 +: 32] = FSM_fft_64_stage_2_0_t412 - FSM_fft_64_stage_2_0_t416;
    FSM_fft_64_stage_2_0_t424 = FSM_fft_64_stage_2_0_t409 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t425 = FSM_fft_64_stage_2_0_t424[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t426 = FSM_fft_64_stage_2_0_t425[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t427 = FSM_fft_64_stage_2_0_t409 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t428 = FSM_fft_64_stage_2_0_t427[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t429 = FSM_fft_64_stage_2_0_t428[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t430 = FSM_fft_64_stage_2_0_t407[FSM_fft_64_stage_2_0_t429 * 32 +: 32];
    FSM_fft_64_stage_2_0_t431 = FSM_fft_64_stage_2_0_t409 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t432 = FSM_fft_64_stage_2_0_t431[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t433 = FSM_fft_64_stage_2_0_t432[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t434 = FSM_fft_64_stage_2_0_t407[FSM_fft_64_stage_2_0_t433 * 32 +: 32];
    FSM_fft_64_stage_2_0_t435 = FSM_fft_64_stage_2_0_t430 + FSM_fft_64_stage_2_0_t434;
    FSM_fft_64_stage_2_0_t436 = FSM_fft_64_stage_2_0_t435[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t437 = FSM_fft_64_stage_2_0_t423;
    FSM_fft_64_stage_2_0_t437[FSM_fft_64_stage_2_0_t426 * 32 +: 32] = FSM_fft_64_stage_2_0_t436;
    FSM_fft_64_stage_2_0_t438 = FSM_fft_64_stage_2_0_t409 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t439 = FSM_fft_64_stage_2_0_t438[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t440 = FSM_fft_64_stage_2_0_t439[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t441 = FSM_fft_64_stage_2_0_t437;
    FSM_fft_64_stage_2_0_t441[FSM_fft_64_stage_2_0_t440 * 32 +: 32] = FSM_fft_64_stage_2_0_t430 - FSM_fft_64_stage_2_0_t434;
    FSM_fft_64_stage_2_0_t442 = 32'b00000000000000000000000000001101 * 32'b00000000000000000000000000000100;
    FSM_fft_64_stage_2_0_t443 = FSM_fft_64_stage_2_0_t442[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t444 = FSM_fft_64_stage_2_0_t443[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t445 = FSM_fft_64_stage_2_0_t443[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t446 = FSM_fft_64_stage_2_0_t441[FSM_fft_64_stage_2_0_t445 * 32 +: 32];
    FSM_fft_64_stage_2_0_t447 = FSM_fft_64_stage_2_0_t443 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t448 = FSM_fft_64_stage_2_0_t447[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t449 = FSM_fft_64_stage_2_0_t448[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t450 = FSM_fft_64_stage_2_0_t441[FSM_fft_64_stage_2_0_t449 * 32 +: 32];
    FSM_fft_64_stage_2_0_t451 = FSM_fft_64_stage_2_0_t446 + FSM_fft_64_stage_2_0_t450;
    FSM_fft_64_stage_2_0_t452 = FSM_fft_64_stage_2_0_t451[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t453 = FSM_fft_64_stage_2_0_t441;
    FSM_fft_64_stage_2_0_t453[FSM_fft_64_stage_2_0_t444 * 32 +: 32] = FSM_fft_64_stage_2_0_t452;
    FSM_fft_64_stage_2_0_t454 = FSM_fft_64_stage_2_0_t443 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t455 = FSM_fft_64_stage_2_0_t454[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t456 = FSM_fft_64_stage_2_0_t455[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t457 = FSM_fft_64_stage_2_0_t453;
    FSM_fft_64_stage_2_0_t457[FSM_fft_64_stage_2_0_t456 * 32 +: 32] = FSM_fft_64_stage_2_0_t446 - FSM_fft_64_stage_2_0_t450;
    FSM_fft_64_stage_2_0_t458 = FSM_fft_64_stage_2_0_t443 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t459 = FSM_fft_64_stage_2_0_t458[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t460 = FSM_fft_64_stage_2_0_t459[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t461 = FSM_fft_64_stage_2_0_t443 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t462 = FSM_fft_64_stage_2_0_t461[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t463 = FSM_fft_64_stage_2_0_t462[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t464 = FSM_fft_64_stage_2_0_t441[FSM_fft_64_stage_2_0_t463 * 32 +: 32];
    FSM_fft_64_stage_2_0_t465 = FSM_fft_64_stage_2_0_t443 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t466 = FSM_fft_64_stage_2_0_t465[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t467 = FSM_fft_64_stage_2_0_t466[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t468 = FSM_fft_64_stage_2_0_t441[FSM_fft_64_stage_2_0_t467 * 32 +: 32];
    FSM_fft_64_stage_2_0_t469 = FSM_fft_64_stage_2_0_t464 + FSM_fft_64_stage_2_0_t468;
    FSM_fft_64_stage_2_0_t470 = FSM_fft_64_stage_2_0_t469[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t471 = FSM_fft_64_stage_2_0_t457;
    FSM_fft_64_stage_2_0_t471[FSM_fft_64_stage_2_0_t460 * 32 +: 32] = FSM_fft_64_stage_2_0_t470;
    FSM_fft_64_stage_2_0_t472 = FSM_fft_64_stage_2_0_t443 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t473 = FSM_fft_64_stage_2_0_t472[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t474 = FSM_fft_64_stage_2_0_t473[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t475 = FSM_fft_64_stage_2_0_t471;
    FSM_fft_64_stage_2_0_t475[FSM_fft_64_stage_2_0_t474 * 32 +: 32] = FSM_fft_64_stage_2_0_t464 - FSM_fft_64_stage_2_0_t468;
    FSM_fft_64_stage_2_0_t476 = 32'b00000000000000000000000000001110 * 32'b00000000000000000000000000000100;
    FSM_fft_64_stage_2_0_t477 = FSM_fft_64_stage_2_0_t476[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t478 = FSM_fft_64_stage_2_0_t477[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t479 = FSM_fft_64_stage_2_0_t477[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t480 = FSM_fft_64_stage_2_0_t475[FSM_fft_64_stage_2_0_t479 * 32 +: 32];
    FSM_fft_64_stage_2_0_t481 = FSM_fft_64_stage_2_0_t477 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t482 = FSM_fft_64_stage_2_0_t481[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t483 = FSM_fft_64_stage_2_0_t482[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t484 = FSM_fft_64_stage_2_0_t475[FSM_fft_64_stage_2_0_t483 * 32 +: 32];
    FSM_fft_64_stage_2_0_t485 = FSM_fft_64_stage_2_0_t480 + FSM_fft_64_stage_2_0_t484;
    FSM_fft_64_stage_2_0_t486 = FSM_fft_64_stage_2_0_t485[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t487 = FSM_fft_64_stage_2_0_t475;
    FSM_fft_64_stage_2_0_t487[FSM_fft_64_stage_2_0_t478 * 32 +: 32] = FSM_fft_64_stage_2_0_t486;
    FSM_fft_64_stage_2_0_t488 = FSM_fft_64_stage_2_0_t477 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t489 = FSM_fft_64_stage_2_0_t488[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t490 = FSM_fft_64_stage_2_0_t489[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t491 = FSM_fft_64_stage_2_0_t487;
    FSM_fft_64_stage_2_0_t491[FSM_fft_64_stage_2_0_t490 * 32 +: 32] = FSM_fft_64_stage_2_0_t480 - FSM_fft_64_stage_2_0_t484;
    FSM_fft_64_stage_2_0_t492 = FSM_fft_64_stage_2_0_t477 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t493 = FSM_fft_64_stage_2_0_t492[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t494 = FSM_fft_64_stage_2_0_t493[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t495 = FSM_fft_64_stage_2_0_t477 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t496 = FSM_fft_64_stage_2_0_t495[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t497 = FSM_fft_64_stage_2_0_t496[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t498 = FSM_fft_64_stage_2_0_t475[FSM_fft_64_stage_2_0_t497 * 32 +: 32];
    FSM_fft_64_stage_2_0_t499 = FSM_fft_64_stage_2_0_t477 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t500 = FSM_fft_64_stage_2_0_t499[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t501 = FSM_fft_64_stage_2_0_t500[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t502 = FSM_fft_64_stage_2_0_t475[FSM_fft_64_stage_2_0_t501 * 32 +: 32];
    FSM_fft_64_stage_2_0_t503 = FSM_fft_64_stage_2_0_t498 + FSM_fft_64_stage_2_0_t502;
    FSM_fft_64_stage_2_0_t504 = FSM_fft_64_stage_2_0_t503[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t505 = FSM_fft_64_stage_2_0_t491;
    FSM_fft_64_stage_2_0_t505[FSM_fft_64_stage_2_0_t494 * 32 +: 32] = FSM_fft_64_stage_2_0_t504;
    FSM_fft_64_stage_2_0_t506 = FSM_fft_64_stage_2_0_t477 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t507 = FSM_fft_64_stage_2_0_t506[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t508 = FSM_fft_64_stage_2_0_t507[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t509 = FSM_fft_64_stage_2_0_t505;
    FSM_fft_64_stage_2_0_t509[FSM_fft_64_stage_2_0_t508 * 32 +: 32] = FSM_fft_64_stage_2_0_t498 - FSM_fft_64_stage_2_0_t502;
    FSM_fft_64_stage_2_0_t510 = 32'b00000000000000000000000000001111 * 32'b00000000000000000000000000000100;
    FSM_fft_64_stage_2_0_t511 = FSM_fft_64_stage_2_0_t510[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t512 = FSM_fft_64_stage_2_0_t511[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t513 = FSM_fft_64_stage_2_0_t511[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t514 = FSM_fft_64_stage_2_0_t509[FSM_fft_64_stage_2_0_t513 * 32 +: 32];
    FSM_fft_64_stage_2_0_t515 = FSM_fft_64_stage_2_0_t511 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t516 = FSM_fft_64_stage_2_0_t515[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t517 = FSM_fft_64_stage_2_0_t516[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t518 = FSM_fft_64_stage_2_0_t509[FSM_fft_64_stage_2_0_t517 * 32 +: 32];
    FSM_fft_64_stage_2_0_t519 = FSM_fft_64_stage_2_0_t514 + FSM_fft_64_stage_2_0_t518;
    FSM_fft_64_stage_2_0_t520 = FSM_fft_64_stage_2_0_t519[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t521 = FSM_fft_64_stage_2_0_t509;
    FSM_fft_64_stage_2_0_t521[FSM_fft_64_stage_2_0_t512 * 32 +: 32] = FSM_fft_64_stage_2_0_t520;
    FSM_fft_64_stage_2_0_t522 = FSM_fft_64_stage_2_0_t511 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t523 = FSM_fft_64_stage_2_0_t522[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t524 = FSM_fft_64_stage_2_0_t523[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t525 = FSM_fft_64_stage_2_0_t521;
    FSM_fft_64_stage_2_0_t525[FSM_fft_64_stage_2_0_t524 * 32 +: 32] = FSM_fft_64_stage_2_0_t514 - FSM_fft_64_stage_2_0_t518;
    FSM_fft_64_stage_2_0_t526 = FSM_fft_64_stage_2_0_t511 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t527 = FSM_fft_64_stage_2_0_t526[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t528 = FSM_fft_64_stage_2_0_t527[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t529 = FSM_fft_64_stage_2_0_t511 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t530 = FSM_fft_64_stage_2_0_t529[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t531 = FSM_fft_64_stage_2_0_t530[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t532 = FSM_fft_64_stage_2_0_t509[FSM_fft_64_stage_2_0_t531 * 32 +: 32];
    FSM_fft_64_stage_2_0_t533 = FSM_fft_64_stage_2_0_t511 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t534 = FSM_fft_64_stage_2_0_t533[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t535 = FSM_fft_64_stage_2_0_t534[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t536 = FSM_fft_64_stage_2_0_t509[FSM_fft_64_stage_2_0_t535 * 32 +: 32];
    FSM_fft_64_stage_2_0_t537 = FSM_fft_64_stage_2_0_t532 + FSM_fft_64_stage_2_0_t536;
    FSM_fft_64_stage_2_0_t538 = FSM_fft_64_stage_2_0_t537[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t539 = FSM_fft_64_stage_2_0_t525;
    FSM_fft_64_stage_2_0_t539[FSM_fft_64_stage_2_0_t528 * 32 +: 32] = FSM_fft_64_stage_2_0_t538;
    FSM_fft_64_stage_2_0_t540 = FSM_fft_64_stage_2_0_t511 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t541 = FSM_fft_64_stage_2_0_t540[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t542 = FSM_fft_64_stage_2_0_t541[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t543 = FSM_fft_64_stage_2_0_t539;
    FSM_fft_64_stage_2_0_t543[FSM_fft_64_stage_2_0_t542 * 32 +: 32] = FSM_fft_64_stage_2_0_t532 - FSM_fft_64_stage_2_0_t536;
    FSM_fft_64_stage_2_0_t544 = FSM_fft_64_stage_2_0_t1[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t545 = FSM_fft_64_stage_2_0_t1[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t546 = i_data_in_imag[FSM_fft_64_stage_2_0_t545 * 32 +: 32];
    FSM_fft_64_stage_2_0_t547 = FSM_fft_64_stage_2_0_t1 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t548 = FSM_fft_64_stage_2_0_t547[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t549 = FSM_fft_64_stage_2_0_t548[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t550 = i_data_in_imag[FSM_fft_64_stage_2_0_t549 * 32 +: 32];
    FSM_fft_64_stage_2_0_t551 = FSM_fft_64_stage_2_0_t546 + FSM_fft_64_stage_2_0_t550;
    FSM_fft_64_stage_2_0_t552 = FSM_fft_64_stage_2_0_t551[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t553 = i_data_in_imag;
    FSM_fft_64_stage_2_0_t553[FSM_fft_64_stage_2_0_t544 * 32 +: 32] = FSM_fft_64_stage_2_0_t552;
    FSM_fft_64_stage_2_0_t554 = FSM_fft_64_stage_2_0_t1 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t555 = FSM_fft_64_stage_2_0_t554[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t556 = FSM_fft_64_stage_2_0_t555[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t557 = FSM_fft_64_stage_2_0_t553;
    FSM_fft_64_stage_2_0_t557[FSM_fft_64_stage_2_0_t556 * 32 +: 32] = FSM_fft_64_stage_2_0_t546 - FSM_fft_64_stage_2_0_t550;
    FSM_fft_64_stage_2_0_t558 = FSM_fft_64_stage_2_0_t1 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t559 = FSM_fft_64_stage_2_0_t558[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t560 = FSM_fft_64_stage_2_0_t559[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t561 = FSM_fft_64_stage_2_0_t1 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t562 = FSM_fft_64_stage_2_0_t561[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t563 = FSM_fft_64_stage_2_0_t562[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t564 = i_data_in_imag[FSM_fft_64_stage_2_0_t563 * 32 +: 32];
    FSM_fft_64_stage_2_0_t565 = FSM_fft_64_stage_2_0_t1 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t566 = FSM_fft_64_stage_2_0_t565[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t567 = FSM_fft_64_stage_2_0_t566[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t568 = i_data_in_imag[FSM_fft_64_stage_2_0_t567 * 32 +: 32];
    FSM_fft_64_stage_2_0_t569 = FSM_fft_64_stage_2_0_t564 + FSM_fft_64_stage_2_0_t568;
    FSM_fft_64_stage_2_0_t570 = FSM_fft_64_stage_2_0_t569[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t571 = FSM_fft_64_stage_2_0_t557;
    FSM_fft_64_stage_2_0_t571[FSM_fft_64_stage_2_0_t560 * 32 +: 32] = FSM_fft_64_stage_2_0_t570;
    FSM_fft_64_stage_2_0_t572 = FSM_fft_64_stage_2_0_t1 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t573 = FSM_fft_64_stage_2_0_t572[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t574 = FSM_fft_64_stage_2_0_t573[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t575 = FSM_fft_64_stage_2_0_t571;
    FSM_fft_64_stage_2_0_t575[FSM_fft_64_stage_2_0_t574 * 32 +: 32] = FSM_fft_64_stage_2_0_t564 - FSM_fft_64_stage_2_0_t568;
    FSM_fft_64_stage_2_0_t576 = FSM_fft_64_stage_2_0_t35[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t577 = FSM_fft_64_stage_2_0_t35[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t578 = FSM_fft_64_stage_2_0_t575[FSM_fft_64_stage_2_0_t577 * 32 +: 32];
    FSM_fft_64_stage_2_0_t579 = FSM_fft_64_stage_2_0_t35 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t580 = FSM_fft_64_stage_2_0_t579[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t581 = FSM_fft_64_stage_2_0_t580[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t582 = FSM_fft_64_stage_2_0_t575[FSM_fft_64_stage_2_0_t581 * 32 +: 32];
    FSM_fft_64_stage_2_0_t583 = FSM_fft_64_stage_2_0_t578 + FSM_fft_64_stage_2_0_t582;
    FSM_fft_64_stage_2_0_t584 = FSM_fft_64_stage_2_0_t583[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t585 = FSM_fft_64_stage_2_0_t575;
    FSM_fft_64_stage_2_0_t585[FSM_fft_64_stage_2_0_t576 * 32 +: 32] = FSM_fft_64_stage_2_0_t584;
    FSM_fft_64_stage_2_0_t586 = FSM_fft_64_stage_2_0_t35 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t587 = FSM_fft_64_stage_2_0_t586[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t588 = FSM_fft_64_stage_2_0_t587[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t589 = FSM_fft_64_stage_2_0_t585;
    FSM_fft_64_stage_2_0_t589[FSM_fft_64_stage_2_0_t588 * 32 +: 32] = FSM_fft_64_stage_2_0_t578 - FSM_fft_64_stage_2_0_t582;
    FSM_fft_64_stage_2_0_t590 = FSM_fft_64_stage_2_0_t35 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t591 = FSM_fft_64_stage_2_0_t590[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t592 = FSM_fft_64_stage_2_0_t591[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t593 = FSM_fft_64_stage_2_0_t35 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t594 = FSM_fft_64_stage_2_0_t593[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t595 = FSM_fft_64_stage_2_0_t594[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t596 = FSM_fft_64_stage_2_0_t575[FSM_fft_64_stage_2_0_t595 * 32 +: 32];
    FSM_fft_64_stage_2_0_t597 = FSM_fft_64_stage_2_0_t35 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t598 = FSM_fft_64_stage_2_0_t597[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t599 = FSM_fft_64_stage_2_0_t598[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t600 = FSM_fft_64_stage_2_0_t575[FSM_fft_64_stage_2_0_t599 * 32 +: 32];
    FSM_fft_64_stage_2_0_t601 = FSM_fft_64_stage_2_0_t596 + FSM_fft_64_stage_2_0_t600;
    FSM_fft_64_stage_2_0_t602 = FSM_fft_64_stage_2_0_t601[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t603 = FSM_fft_64_stage_2_0_t589;
    FSM_fft_64_stage_2_0_t603[FSM_fft_64_stage_2_0_t592 * 32 +: 32] = FSM_fft_64_stage_2_0_t602;
    FSM_fft_64_stage_2_0_t604 = FSM_fft_64_stage_2_0_t35 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t605 = FSM_fft_64_stage_2_0_t604[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t606 = FSM_fft_64_stage_2_0_t605[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t607 = FSM_fft_64_stage_2_0_t603;
    FSM_fft_64_stage_2_0_t607[FSM_fft_64_stage_2_0_t606 * 32 +: 32] = FSM_fft_64_stage_2_0_t596 - FSM_fft_64_stage_2_0_t600;
    FSM_fft_64_stage_2_0_t608 = FSM_fft_64_stage_2_0_t69[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t609 = FSM_fft_64_stage_2_0_t69[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t610 = FSM_fft_64_stage_2_0_t607[FSM_fft_64_stage_2_0_t609 * 32 +: 32];
    FSM_fft_64_stage_2_0_t611 = FSM_fft_64_stage_2_0_t69 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t612 = FSM_fft_64_stage_2_0_t611[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t613 = FSM_fft_64_stage_2_0_t612[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t614 = FSM_fft_64_stage_2_0_t607[FSM_fft_64_stage_2_0_t613 * 32 +: 32];
    FSM_fft_64_stage_2_0_t615 = FSM_fft_64_stage_2_0_t610 + FSM_fft_64_stage_2_0_t614;
    FSM_fft_64_stage_2_0_t616 = FSM_fft_64_stage_2_0_t615[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t617 = FSM_fft_64_stage_2_0_t607;
    FSM_fft_64_stage_2_0_t617[FSM_fft_64_stage_2_0_t608 * 32 +: 32] = FSM_fft_64_stage_2_0_t616;
    FSM_fft_64_stage_2_0_t618 = FSM_fft_64_stage_2_0_t69 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t619 = FSM_fft_64_stage_2_0_t618[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t620 = FSM_fft_64_stage_2_0_t619[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t621 = FSM_fft_64_stage_2_0_t617;
    FSM_fft_64_stage_2_0_t621[FSM_fft_64_stage_2_0_t620 * 32 +: 32] = FSM_fft_64_stage_2_0_t610 - FSM_fft_64_stage_2_0_t614;
    FSM_fft_64_stage_2_0_t622 = FSM_fft_64_stage_2_0_t69 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t623 = FSM_fft_64_stage_2_0_t622[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t624 = FSM_fft_64_stage_2_0_t623[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t625 = FSM_fft_64_stage_2_0_t69 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t626 = FSM_fft_64_stage_2_0_t625[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t627 = FSM_fft_64_stage_2_0_t626[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t628 = FSM_fft_64_stage_2_0_t607[FSM_fft_64_stage_2_0_t627 * 32 +: 32];
    FSM_fft_64_stage_2_0_t629 = FSM_fft_64_stage_2_0_t69 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t630 = FSM_fft_64_stage_2_0_t629[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t631 = FSM_fft_64_stage_2_0_t630[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t632 = FSM_fft_64_stage_2_0_t607[FSM_fft_64_stage_2_0_t631 * 32 +: 32];
    FSM_fft_64_stage_2_0_t633 = FSM_fft_64_stage_2_0_t628 + FSM_fft_64_stage_2_0_t632;
    FSM_fft_64_stage_2_0_t634 = FSM_fft_64_stage_2_0_t633[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t635 = FSM_fft_64_stage_2_0_t621;
    FSM_fft_64_stage_2_0_t635[FSM_fft_64_stage_2_0_t624 * 32 +: 32] = FSM_fft_64_stage_2_0_t634;
    FSM_fft_64_stage_2_0_t636 = FSM_fft_64_stage_2_0_t69 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t637 = FSM_fft_64_stage_2_0_t636[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t638 = FSM_fft_64_stage_2_0_t637[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t639 = FSM_fft_64_stage_2_0_t635;
    FSM_fft_64_stage_2_0_t639[FSM_fft_64_stage_2_0_t638 * 32 +: 32] = FSM_fft_64_stage_2_0_t628 - FSM_fft_64_stage_2_0_t632;
    FSM_fft_64_stage_2_0_t640 = FSM_fft_64_stage_2_0_t103[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t641 = FSM_fft_64_stage_2_0_t103[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t642 = FSM_fft_64_stage_2_0_t639[FSM_fft_64_stage_2_0_t641 * 32 +: 32];
    FSM_fft_64_stage_2_0_t643 = FSM_fft_64_stage_2_0_t103 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t644 = FSM_fft_64_stage_2_0_t643[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t645 = FSM_fft_64_stage_2_0_t644[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t646 = FSM_fft_64_stage_2_0_t639[FSM_fft_64_stage_2_0_t645 * 32 +: 32];
    FSM_fft_64_stage_2_0_t647 = FSM_fft_64_stage_2_0_t642 + FSM_fft_64_stage_2_0_t646;
    FSM_fft_64_stage_2_0_t648 = FSM_fft_64_stage_2_0_t647[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t649 = FSM_fft_64_stage_2_0_t639;
    FSM_fft_64_stage_2_0_t649[FSM_fft_64_stage_2_0_t640 * 32 +: 32] = FSM_fft_64_stage_2_0_t648;
    FSM_fft_64_stage_2_0_t650 = FSM_fft_64_stage_2_0_t103 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t651 = FSM_fft_64_stage_2_0_t650[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t652 = FSM_fft_64_stage_2_0_t651[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t653 = FSM_fft_64_stage_2_0_t649;
    FSM_fft_64_stage_2_0_t653[FSM_fft_64_stage_2_0_t652 * 32 +: 32] = FSM_fft_64_stage_2_0_t642 - FSM_fft_64_stage_2_0_t646;
    FSM_fft_64_stage_2_0_t654 = FSM_fft_64_stage_2_0_t103 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t655 = FSM_fft_64_stage_2_0_t654[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t656 = FSM_fft_64_stage_2_0_t655[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t657 = FSM_fft_64_stage_2_0_t103 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t658 = FSM_fft_64_stage_2_0_t657[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t659 = FSM_fft_64_stage_2_0_t658[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t660 = FSM_fft_64_stage_2_0_t639[FSM_fft_64_stage_2_0_t659 * 32 +: 32];
    FSM_fft_64_stage_2_0_t661 = FSM_fft_64_stage_2_0_t103 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t662 = FSM_fft_64_stage_2_0_t661[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t663 = FSM_fft_64_stage_2_0_t662[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t664 = FSM_fft_64_stage_2_0_t639[FSM_fft_64_stage_2_0_t663 * 32 +: 32];
    FSM_fft_64_stage_2_0_t665 = FSM_fft_64_stage_2_0_t660 + FSM_fft_64_stage_2_0_t664;
    FSM_fft_64_stage_2_0_t666 = FSM_fft_64_stage_2_0_t665[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t667 = FSM_fft_64_stage_2_0_t653;
    FSM_fft_64_stage_2_0_t667[FSM_fft_64_stage_2_0_t656 * 32 +: 32] = FSM_fft_64_stage_2_0_t666;
    FSM_fft_64_stage_2_0_t668 = FSM_fft_64_stage_2_0_t103 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t669 = FSM_fft_64_stage_2_0_t668[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t670 = FSM_fft_64_stage_2_0_t669[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t671 = FSM_fft_64_stage_2_0_t667;
    FSM_fft_64_stage_2_0_t671[FSM_fft_64_stage_2_0_t670 * 32 +: 32] = FSM_fft_64_stage_2_0_t660 - FSM_fft_64_stage_2_0_t664;
    FSM_fft_64_stage_2_0_t672 = FSM_fft_64_stage_2_0_t137[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t673 = FSM_fft_64_stage_2_0_t137[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t674 = FSM_fft_64_stage_2_0_t671[FSM_fft_64_stage_2_0_t673 * 32 +: 32];
    FSM_fft_64_stage_2_0_t675 = FSM_fft_64_stage_2_0_t137 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t676 = FSM_fft_64_stage_2_0_t675[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t677 = FSM_fft_64_stage_2_0_t676[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t678 = FSM_fft_64_stage_2_0_t671[FSM_fft_64_stage_2_0_t677 * 32 +: 32];
    FSM_fft_64_stage_2_0_t679 = FSM_fft_64_stage_2_0_t674 + FSM_fft_64_stage_2_0_t678;
    FSM_fft_64_stage_2_0_t680 = FSM_fft_64_stage_2_0_t679[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t681 = FSM_fft_64_stage_2_0_t671;
    FSM_fft_64_stage_2_0_t681[FSM_fft_64_stage_2_0_t672 * 32 +: 32] = FSM_fft_64_stage_2_0_t680;
    FSM_fft_64_stage_2_0_t682 = FSM_fft_64_stage_2_0_t137 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t683 = FSM_fft_64_stage_2_0_t682[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t684 = FSM_fft_64_stage_2_0_t683[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t685 = FSM_fft_64_stage_2_0_t681;
    FSM_fft_64_stage_2_0_t685[FSM_fft_64_stage_2_0_t684 * 32 +: 32] = FSM_fft_64_stage_2_0_t674 - FSM_fft_64_stage_2_0_t678;
    FSM_fft_64_stage_2_0_t686 = FSM_fft_64_stage_2_0_t137 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t687 = FSM_fft_64_stage_2_0_t686[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t688 = FSM_fft_64_stage_2_0_t687[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t689 = FSM_fft_64_stage_2_0_t137 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t690 = FSM_fft_64_stage_2_0_t689[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t691 = FSM_fft_64_stage_2_0_t690[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t692 = FSM_fft_64_stage_2_0_t671[FSM_fft_64_stage_2_0_t691 * 32 +: 32];
    FSM_fft_64_stage_2_0_t693 = FSM_fft_64_stage_2_0_t137 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t694 = FSM_fft_64_stage_2_0_t693[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t695 = FSM_fft_64_stage_2_0_t694[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t696 = FSM_fft_64_stage_2_0_t671[FSM_fft_64_stage_2_0_t695 * 32 +: 32];
    FSM_fft_64_stage_2_0_t697 = FSM_fft_64_stage_2_0_t692 + FSM_fft_64_stage_2_0_t696;
    FSM_fft_64_stage_2_0_t698 = FSM_fft_64_stage_2_0_t697[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t699 = FSM_fft_64_stage_2_0_t685;
    FSM_fft_64_stage_2_0_t699[FSM_fft_64_stage_2_0_t688 * 32 +: 32] = FSM_fft_64_stage_2_0_t698;
    FSM_fft_64_stage_2_0_t700 = FSM_fft_64_stage_2_0_t137 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t701 = FSM_fft_64_stage_2_0_t700[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t702 = FSM_fft_64_stage_2_0_t701[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t703 = FSM_fft_64_stage_2_0_t699;
    FSM_fft_64_stage_2_0_t703[FSM_fft_64_stage_2_0_t702 * 32 +: 32] = FSM_fft_64_stage_2_0_t692 - FSM_fft_64_stage_2_0_t696;
    FSM_fft_64_stage_2_0_t704 = FSM_fft_64_stage_2_0_t171[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t705 = FSM_fft_64_stage_2_0_t171[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t706 = FSM_fft_64_stage_2_0_t703[FSM_fft_64_stage_2_0_t705 * 32 +: 32];
    FSM_fft_64_stage_2_0_t707 = FSM_fft_64_stage_2_0_t171 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t708 = FSM_fft_64_stage_2_0_t707[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t709 = FSM_fft_64_stage_2_0_t708[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t710 = FSM_fft_64_stage_2_0_t703[FSM_fft_64_stage_2_0_t709 * 32 +: 32];
    FSM_fft_64_stage_2_0_t711 = FSM_fft_64_stage_2_0_t706 + FSM_fft_64_stage_2_0_t710;
    FSM_fft_64_stage_2_0_t712 = FSM_fft_64_stage_2_0_t711[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t713 = FSM_fft_64_stage_2_0_t703;
    FSM_fft_64_stage_2_0_t713[FSM_fft_64_stage_2_0_t704 * 32 +: 32] = FSM_fft_64_stage_2_0_t712;
    FSM_fft_64_stage_2_0_t714 = FSM_fft_64_stage_2_0_t171 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t715 = FSM_fft_64_stage_2_0_t714[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t716 = FSM_fft_64_stage_2_0_t715[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t717 = FSM_fft_64_stage_2_0_t713;
    FSM_fft_64_stage_2_0_t717[FSM_fft_64_stage_2_0_t716 * 32 +: 32] = FSM_fft_64_stage_2_0_t706 - FSM_fft_64_stage_2_0_t710;
    FSM_fft_64_stage_2_0_t718 = FSM_fft_64_stage_2_0_t171 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t719 = FSM_fft_64_stage_2_0_t718[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t720 = FSM_fft_64_stage_2_0_t719[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t721 = FSM_fft_64_stage_2_0_t171 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t722 = FSM_fft_64_stage_2_0_t721[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t723 = FSM_fft_64_stage_2_0_t722[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t724 = FSM_fft_64_stage_2_0_t703[FSM_fft_64_stage_2_0_t723 * 32 +: 32];
    FSM_fft_64_stage_2_0_t725 = FSM_fft_64_stage_2_0_t171 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t726 = FSM_fft_64_stage_2_0_t725[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t727 = FSM_fft_64_stage_2_0_t726[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t728 = FSM_fft_64_stage_2_0_t703[FSM_fft_64_stage_2_0_t727 * 32 +: 32];
    FSM_fft_64_stage_2_0_t729 = FSM_fft_64_stage_2_0_t724 + FSM_fft_64_stage_2_0_t728;
    FSM_fft_64_stage_2_0_t730 = FSM_fft_64_stage_2_0_t729[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t731 = FSM_fft_64_stage_2_0_t717;
    FSM_fft_64_stage_2_0_t731[FSM_fft_64_stage_2_0_t720 * 32 +: 32] = FSM_fft_64_stage_2_0_t730;
    FSM_fft_64_stage_2_0_t732 = FSM_fft_64_stage_2_0_t171 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t733 = FSM_fft_64_stage_2_0_t732[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t734 = FSM_fft_64_stage_2_0_t733[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t735 = FSM_fft_64_stage_2_0_t731;
    FSM_fft_64_stage_2_0_t735[FSM_fft_64_stage_2_0_t734 * 32 +: 32] = FSM_fft_64_stage_2_0_t724 - FSM_fft_64_stage_2_0_t728;
    FSM_fft_64_stage_2_0_t736 = FSM_fft_64_stage_2_0_t205[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t737 = FSM_fft_64_stage_2_0_t205[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t738 = FSM_fft_64_stage_2_0_t735[FSM_fft_64_stage_2_0_t737 * 32 +: 32];
    FSM_fft_64_stage_2_0_t739 = FSM_fft_64_stage_2_0_t205 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t740 = FSM_fft_64_stage_2_0_t739[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t741 = FSM_fft_64_stage_2_0_t740[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t742 = FSM_fft_64_stage_2_0_t735[FSM_fft_64_stage_2_0_t741 * 32 +: 32];
    FSM_fft_64_stage_2_0_t743 = FSM_fft_64_stage_2_0_t738 + FSM_fft_64_stage_2_0_t742;
    FSM_fft_64_stage_2_0_t744 = FSM_fft_64_stage_2_0_t743[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t745 = FSM_fft_64_stage_2_0_t735;
    FSM_fft_64_stage_2_0_t745[FSM_fft_64_stage_2_0_t736 * 32 +: 32] = FSM_fft_64_stage_2_0_t744;
    FSM_fft_64_stage_2_0_t746 = FSM_fft_64_stage_2_0_t205 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t747 = FSM_fft_64_stage_2_0_t746[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t748 = FSM_fft_64_stage_2_0_t747[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t749 = FSM_fft_64_stage_2_0_t745;
    FSM_fft_64_stage_2_0_t749[FSM_fft_64_stage_2_0_t748 * 32 +: 32] = FSM_fft_64_stage_2_0_t738 - FSM_fft_64_stage_2_0_t742;
    FSM_fft_64_stage_2_0_t750 = FSM_fft_64_stage_2_0_t205 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t751 = FSM_fft_64_stage_2_0_t750[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t752 = FSM_fft_64_stage_2_0_t751[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t753 = FSM_fft_64_stage_2_0_t205 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t754 = FSM_fft_64_stage_2_0_t753[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t755 = FSM_fft_64_stage_2_0_t754[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t756 = FSM_fft_64_stage_2_0_t735[FSM_fft_64_stage_2_0_t755 * 32 +: 32];
    FSM_fft_64_stage_2_0_t757 = FSM_fft_64_stage_2_0_t205 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t758 = FSM_fft_64_stage_2_0_t757[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t759 = FSM_fft_64_stage_2_0_t758[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t760 = FSM_fft_64_stage_2_0_t735[FSM_fft_64_stage_2_0_t759 * 32 +: 32];
    FSM_fft_64_stage_2_0_t761 = FSM_fft_64_stage_2_0_t756 + FSM_fft_64_stage_2_0_t760;
    FSM_fft_64_stage_2_0_t762 = FSM_fft_64_stage_2_0_t761[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t763 = FSM_fft_64_stage_2_0_t749;
    FSM_fft_64_stage_2_0_t763[FSM_fft_64_stage_2_0_t752 * 32 +: 32] = FSM_fft_64_stage_2_0_t762;
    FSM_fft_64_stage_2_0_t764 = FSM_fft_64_stage_2_0_t205 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t765 = FSM_fft_64_stage_2_0_t764[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t766 = FSM_fft_64_stage_2_0_t765[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t767 = FSM_fft_64_stage_2_0_t763;
    FSM_fft_64_stage_2_0_t767[FSM_fft_64_stage_2_0_t766 * 32 +: 32] = FSM_fft_64_stage_2_0_t756 - FSM_fft_64_stage_2_0_t760;
    FSM_fft_64_stage_2_0_t768 = FSM_fft_64_stage_2_0_t239[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t769 = FSM_fft_64_stage_2_0_t239[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t770 = FSM_fft_64_stage_2_0_t767[FSM_fft_64_stage_2_0_t769 * 32 +: 32];
    FSM_fft_64_stage_2_0_t771 = FSM_fft_64_stage_2_0_t239 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t772 = FSM_fft_64_stage_2_0_t771[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t773 = FSM_fft_64_stage_2_0_t772[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t774 = FSM_fft_64_stage_2_0_t767[FSM_fft_64_stage_2_0_t773 * 32 +: 32];
    FSM_fft_64_stage_2_0_t775 = FSM_fft_64_stage_2_0_t770 + FSM_fft_64_stage_2_0_t774;
    FSM_fft_64_stage_2_0_t776 = FSM_fft_64_stage_2_0_t775[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t777 = FSM_fft_64_stage_2_0_t767;
    FSM_fft_64_stage_2_0_t777[FSM_fft_64_stage_2_0_t768 * 32 +: 32] = FSM_fft_64_stage_2_0_t776;
    FSM_fft_64_stage_2_0_t778 = FSM_fft_64_stage_2_0_t239 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t779 = FSM_fft_64_stage_2_0_t778[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t780 = FSM_fft_64_stage_2_0_t779[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t781 = FSM_fft_64_stage_2_0_t777;
    FSM_fft_64_stage_2_0_t781[FSM_fft_64_stage_2_0_t780 * 32 +: 32] = FSM_fft_64_stage_2_0_t770 - FSM_fft_64_stage_2_0_t774;
    FSM_fft_64_stage_2_0_t782 = FSM_fft_64_stage_2_0_t239 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t783 = FSM_fft_64_stage_2_0_t782[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t784 = FSM_fft_64_stage_2_0_t783[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t785 = FSM_fft_64_stage_2_0_t239 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t786 = FSM_fft_64_stage_2_0_t785[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t787 = FSM_fft_64_stage_2_0_t786[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t788 = FSM_fft_64_stage_2_0_t767[FSM_fft_64_stage_2_0_t787 * 32 +: 32];
    FSM_fft_64_stage_2_0_t789 = FSM_fft_64_stage_2_0_t239 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t790 = FSM_fft_64_stage_2_0_t789[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t791 = FSM_fft_64_stage_2_0_t790[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t792 = FSM_fft_64_stage_2_0_t767[FSM_fft_64_stage_2_0_t791 * 32 +: 32];
    FSM_fft_64_stage_2_0_t793 = FSM_fft_64_stage_2_0_t788 + FSM_fft_64_stage_2_0_t792;
    FSM_fft_64_stage_2_0_t794 = FSM_fft_64_stage_2_0_t793[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t795 = FSM_fft_64_stage_2_0_t781;
    FSM_fft_64_stage_2_0_t795[FSM_fft_64_stage_2_0_t784 * 32 +: 32] = FSM_fft_64_stage_2_0_t794;
    FSM_fft_64_stage_2_0_t796 = FSM_fft_64_stage_2_0_t239 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t797 = FSM_fft_64_stage_2_0_t796[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t798 = FSM_fft_64_stage_2_0_t797[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t799 = FSM_fft_64_stage_2_0_t795;
    FSM_fft_64_stage_2_0_t799[FSM_fft_64_stage_2_0_t798 * 32 +: 32] = FSM_fft_64_stage_2_0_t788 - FSM_fft_64_stage_2_0_t792;
    FSM_fft_64_stage_2_0_t800 = FSM_fft_64_stage_2_0_t273[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t801 = FSM_fft_64_stage_2_0_t273[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t802 = FSM_fft_64_stage_2_0_t799[FSM_fft_64_stage_2_0_t801 * 32 +: 32];
    FSM_fft_64_stage_2_0_t803 = FSM_fft_64_stage_2_0_t273 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t804 = FSM_fft_64_stage_2_0_t803[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t805 = FSM_fft_64_stage_2_0_t804[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t806 = FSM_fft_64_stage_2_0_t799[FSM_fft_64_stage_2_0_t805 * 32 +: 32];
    FSM_fft_64_stage_2_0_t807 = FSM_fft_64_stage_2_0_t802 + FSM_fft_64_stage_2_0_t806;
    FSM_fft_64_stage_2_0_t808 = FSM_fft_64_stage_2_0_t807[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t809 = FSM_fft_64_stage_2_0_t799;
    FSM_fft_64_stage_2_0_t809[FSM_fft_64_stage_2_0_t800 * 32 +: 32] = FSM_fft_64_stage_2_0_t808;
    FSM_fft_64_stage_2_0_t810 = FSM_fft_64_stage_2_0_t273 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t811 = FSM_fft_64_stage_2_0_t810[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t812 = FSM_fft_64_stage_2_0_t811[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t813 = FSM_fft_64_stage_2_0_t809;
    FSM_fft_64_stage_2_0_t813[FSM_fft_64_stage_2_0_t812 * 32 +: 32] = FSM_fft_64_stage_2_0_t802 - FSM_fft_64_stage_2_0_t806;
    FSM_fft_64_stage_2_0_t814 = FSM_fft_64_stage_2_0_t273 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t815 = FSM_fft_64_stage_2_0_t814[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t816 = FSM_fft_64_stage_2_0_t815[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t817 = FSM_fft_64_stage_2_0_t273 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t818 = FSM_fft_64_stage_2_0_t817[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t819 = FSM_fft_64_stage_2_0_t818[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t820 = FSM_fft_64_stage_2_0_t799[FSM_fft_64_stage_2_0_t819 * 32 +: 32];
    FSM_fft_64_stage_2_0_t821 = FSM_fft_64_stage_2_0_t273 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t822 = FSM_fft_64_stage_2_0_t821[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t823 = FSM_fft_64_stage_2_0_t822[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t824 = FSM_fft_64_stage_2_0_t799[FSM_fft_64_stage_2_0_t823 * 32 +: 32];
    FSM_fft_64_stage_2_0_t825 = FSM_fft_64_stage_2_0_t820 + FSM_fft_64_stage_2_0_t824;
    FSM_fft_64_stage_2_0_t826 = FSM_fft_64_stage_2_0_t825[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t827 = FSM_fft_64_stage_2_0_t813;
    FSM_fft_64_stage_2_0_t827[FSM_fft_64_stage_2_0_t816 * 32 +: 32] = FSM_fft_64_stage_2_0_t826;
    FSM_fft_64_stage_2_0_t828 = FSM_fft_64_stage_2_0_t273 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t829 = FSM_fft_64_stage_2_0_t828[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t830 = FSM_fft_64_stage_2_0_t829[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t831 = FSM_fft_64_stage_2_0_t827;
    FSM_fft_64_stage_2_0_t831[FSM_fft_64_stage_2_0_t830 * 32 +: 32] = FSM_fft_64_stage_2_0_t820 - FSM_fft_64_stage_2_0_t824;
    FSM_fft_64_stage_2_0_t832 = FSM_fft_64_stage_2_0_t307[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t833 = FSM_fft_64_stage_2_0_t307[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t834 = FSM_fft_64_stage_2_0_t831[FSM_fft_64_stage_2_0_t833 * 32 +: 32];
    FSM_fft_64_stage_2_0_t835 = FSM_fft_64_stage_2_0_t307 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t836 = FSM_fft_64_stage_2_0_t835[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t837 = FSM_fft_64_stage_2_0_t836[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t838 = FSM_fft_64_stage_2_0_t831[FSM_fft_64_stage_2_0_t837 * 32 +: 32];
    FSM_fft_64_stage_2_0_t839 = FSM_fft_64_stage_2_0_t834 + FSM_fft_64_stage_2_0_t838;
    FSM_fft_64_stage_2_0_t840 = FSM_fft_64_stage_2_0_t839[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t841 = FSM_fft_64_stage_2_0_t831;
    FSM_fft_64_stage_2_0_t841[FSM_fft_64_stage_2_0_t832 * 32 +: 32] = FSM_fft_64_stage_2_0_t840;
    FSM_fft_64_stage_2_0_t842 = FSM_fft_64_stage_2_0_t307 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t843 = FSM_fft_64_stage_2_0_t842[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t844 = FSM_fft_64_stage_2_0_t843[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t845 = FSM_fft_64_stage_2_0_t841;
    FSM_fft_64_stage_2_0_t845[FSM_fft_64_stage_2_0_t844 * 32 +: 32] = FSM_fft_64_stage_2_0_t834 - FSM_fft_64_stage_2_0_t838;
    FSM_fft_64_stage_2_0_t846 = FSM_fft_64_stage_2_0_t307 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t847 = FSM_fft_64_stage_2_0_t846[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t848 = FSM_fft_64_stage_2_0_t847[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t849 = FSM_fft_64_stage_2_0_t307 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t850 = FSM_fft_64_stage_2_0_t849[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t851 = FSM_fft_64_stage_2_0_t850[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t852 = FSM_fft_64_stage_2_0_t831[FSM_fft_64_stage_2_0_t851 * 32 +: 32];
    FSM_fft_64_stage_2_0_t853 = FSM_fft_64_stage_2_0_t307 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t854 = FSM_fft_64_stage_2_0_t853[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t855 = FSM_fft_64_stage_2_0_t854[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t856 = FSM_fft_64_stage_2_0_t831[FSM_fft_64_stage_2_0_t855 * 32 +: 32];
    FSM_fft_64_stage_2_0_t857 = FSM_fft_64_stage_2_0_t852 + FSM_fft_64_stage_2_0_t856;
    FSM_fft_64_stage_2_0_t858 = FSM_fft_64_stage_2_0_t857[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t859 = FSM_fft_64_stage_2_0_t845;
    FSM_fft_64_stage_2_0_t859[FSM_fft_64_stage_2_0_t848 * 32 +: 32] = FSM_fft_64_stage_2_0_t858;
    FSM_fft_64_stage_2_0_t860 = FSM_fft_64_stage_2_0_t307 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t861 = FSM_fft_64_stage_2_0_t860[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t862 = FSM_fft_64_stage_2_0_t861[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t863 = FSM_fft_64_stage_2_0_t859;
    FSM_fft_64_stage_2_0_t863[FSM_fft_64_stage_2_0_t862 * 32 +: 32] = FSM_fft_64_stage_2_0_t852 - FSM_fft_64_stage_2_0_t856;
    FSM_fft_64_stage_2_0_t864 = FSM_fft_64_stage_2_0_t341[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t865 = FSM_fft_64_stage_2_0_t341[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t866 = FSM_fft_64_stage_2_0_t863[FSM_fft_64_stage_2_0_t865 * 32 +: 32];
    FSM_fft_64_stage_2_0_t867 = FSM_fft_64_stage_2_0_t341 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t868 = FSM_fft_64_stage_2_0_t867[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t869 = FSM_fft_64_stage_2_0_t868[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t870 = FSM_fft_64_stage_2_0_t863[FSM_fft_64_stage_2_0_t869 * 32 +: 32];
    FSM_fft_64_stage_2_0_t871 = FSM_fft_64_stage_2_0_t866 + FSM_fft_64_stage_2_0_t870;
    FSM_fft_64_stage_2_0_t872 = FSM_fft_64_stage_2_0_t871[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t873 = FSM_fft_64_stage_2_0_t863;
    FSM_fft_64_stage_2_0_t873[FSM_fft_64_stage_2_0_t864 * 32 +: 32] = FSM_fft_64_stage_2_0_t872;
    FSM_fft_64_stage_2_0_t874 = FSM_fft_64_stage_2_0_t341 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t875 = FSM_fft_64_stage_2_0_t874[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t876 = FSM_fft_64_stage_2_0_t875[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t877 = FSM_fft_64_stage_2_0_t873;
    FSM_fft_64_stage_2_0_t877[FSM_fft_64_stage_2_0_t876 * 32 +: 32] = FSM_fft_64_stage_2_0_t866 - FSM_fft_64_stage_2_0_t870;
    FSM_fft_64_stage_2_0_t878 = FSM_fft_64_stage_2_0_t341 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t879 = FSM_fft_64_stage_2_0_t878[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t880 = FSM_fft_64_stage_2_0_t879[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t881 = FSM_fft_64_stage_2_0_t341 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t882 = FSM_fft_64_stage_2_0_t881[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t883 = FSM_fft_64_stage_2_0_t882[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t884 = FSM_fft_64_stage_2_0_t863[FSM_fft_64_stage_2_0_t883 * 32 +: 32];
    FSM_fft_64_stage_2_0_t885 = FSM_fft_64_stage_2_0_t341 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t886 = FSM_fft_64_stage_2_0_t885[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t887 = FSM_fft_64_stage_2_0_t886[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t888 = FSM_fft_64_stage_2_0_t863[FSM_fft_64_stage_2_0_t887 * 32 +: 32];
    FSM_fft_64_stage_2_0_t889 = FSM_fft_64_stage_2_0_t884 + FSM_fft_64_stage_2_0_t888;
    FSM_fft_64_stage_2_0_t890 = FSM_fft_64_stage_2_0_t889[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t891 = FSM_fft_64_stage_2_0_t877;
    FSM_fft_64_stage_2_0_t891[FSM_fft_64_stage_2_0_t880 * 32 +: 32] = FSM_fft_64_stage_2_0_t890;
    FSM_fft_64_stage_2_0_t892 = FSM_fft_64_stage_2_0_t341 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t893 = FSM_fft_64_stage_2_0_t892[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t894 = FSM_fft_64_stage_2_0_t893[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t895 = FSM_fft_64_stage_2_0_t891;
    FSM_fft_64_stage_2_0_t895[FSM_fft_64_stage_2_0_t894 * 32 +: 32] = FSM_fft_64_stage_2_0_t884 - FSM_fft_64_stage_2_0_t888;
    FSM_fft_64_stage_2_0_t896 = FSM_fft_64_stage_2_0_t375[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t897 = FSM_fft_64_stage_2_0_t375[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t898 = FSM_fft_64_stage_2_0_t895[FSM_fft_64_stage_2_0_t897 * 32 +: 32];
    FSM_fft_64_stage_2_0_t899 = FSM_fft_64_stage_2_0_t375 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t900 = FSM_fft_64_stage_2_0_t899[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t901 = FSM_fft_64_stage_2_0_t900[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t902 = FSM_fft_64_stage_2_0_t895[FSM_fft_64_stage_2_0_t901 * 32 +: 32];
    FSM_fft_64_stage_2_0_t903 = FSM_fft_64_stage_2_0_t898 + FSM_fft_64_stage_2_0_t902;
    FSM_fft_64_stage_2_0_t904 = FSM_fft_64_stage_2_0_t903[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t905 = FSM_fft_64_stage_2_0_t895;
    FSM_fft_64_stage_2_0_t905[FSM_fft_64_stage_2_0_t896 * 32 +: 32] = FSM_fft_64_stage_2_0_t904;
    FSM_fft_64_stage_2_0_t906 = FSM_fft_64_stage_2_0_t375 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t907 = FSM_fft_64_stage_2_0_t906[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t908 = FSM_fft_64_stage_2_0_t907[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t909 = FSM_fft_64_stage_2_0_t905;
    FSM_fft_64_stage_2_0_t909[FSM_fft_64_stage_2_0_t908 * 32 +: 32] = FSM_fft_64_stage_2_0_t898 - FSM_fft_64_stage_2_0_t902;
    FSM_fft_64_stage_2_0_t910 = FSM_fft_64_stage_2_0_t375 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t911 = FSM_fft_64_stage_2_0_t910[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t912 = FSM_fft_64_stage_2_0_t911[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t913 = FSM_fft_64_stage_2_0_t375 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t914 = FSM_fft_64_stage_2_0_t913[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t915 = FSM_fft_64_stage_2_0_t914[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t916 = FSM_fft_64_stage_2_0_t895[FSM_fft_64_stage_2_0_t915 * 32 +: 32];
    FSM_fft_64_stage_2_0_t917 = FSM_fft_64_stage_2_0_t375 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t918 = FSM_fft_64_stage_2_0_t917[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t919 = FSM_fft_64_stage_2_0_t918[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t920 = FSM_fft_64_stage_2_0_t895[FSM_fft_64_stage_2_0_t919 * 32 +: 32];
    FSM_fft_64_stage_2_0_t921 = FSM_fft_64_stage_2_0_t916 + FSM_fft_64_stage_2_0_t920;
    FSM_fft_64_stage_2_0_t922 = FSM_fft_64_stage_2_0_t921[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t923 = FSM_fft_64_stage_2_0_t909;
    FSM_fft_64_stage_2_0_t923[FSM_fft_64_stage_2_0_t912 * 32 +: 32] = FSM_fft_64_stage_2_0_t922;
    FSM_fft_64_stage_2_0_t924 = FSM_fft_64_stage_2_0_t375 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t925 = FSM_fft_64_stage_2_0_t924[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t926 = FSM_fft_64_stage_2_0_t925[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t927 = FSM_fft_64_stage_2_0_t923;
    FSM_fft_64_stage_2_0_t927[FSM_fft_64_stage_2_0_t926 * 32 +: 32] = FSM_fft_64_stage_2_0_t916 - FSM_fft_64_stage_2_0_t920;
    FSM_fft_64_stage_2_0_t928 = FSM_fft_64_stage_2_0_t409[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t929 = FSM_fft_64_stage_2_0_t409[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t930 = FSM_fft_64_stage_2_0_t927[FSM_fft_64_stage_2_0_t929 * 32 +: 32];
    FSM_fft_64_stage_2_0_t931 = FSM_fft_64_stage_2_0_t409 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t932 = FSM_fft_64_stage_2_0_t931[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t933 = FSM_fft_64_stage_2_0_t932[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t934 = FSM_fft_64_stage_2_0_t927[FSM_fft_64_stage_2_0_t933 * 32 +: 32];
    FSM_fft_64_stage_2_0_t935 = FSM_fft_64_stage_2_0_t930 + FSM_fft_64_stage_2_0_t934;
    FSM_fft_64_stage_2_0_t936 = FSM_fft_64_stage_2_0_t935[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t937 = FSM_fft_64_stage_2_0_t927;
    FSM_fft_64_stage_2_0_t937[FSM_fft_64_stage_2_0_t928 * 32 +: 32] = FSM_fft_64_stage_2_0_t936;
    FSM_fft_64_stage_2_0_t938 = FSM_fft_64_stage_2_0_t409 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t939 = FSM_fft_64_stage_2_0_t938[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t940 = FSM_fft_64_stage_2_0_t939[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t941 = FSM_fft_64_stage_2_0_t937;
    FSM_fft_64_stage_2_0_t941[FSM_fft_64_stage_2_0_t940 * 32 +: 32] = FSM_fft_64_stage_2_0_t930 - FSM_fft_64_stage_2_0_t934;
    FSM_fft_64_stage_2_0_t942 = FSM_fft_64_stage_2_0_t409 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t943 = FSM_fft_64_stage_2_0_t942[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t944 = FSM_fft_64_stage_2_0_t943[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t945 = FSM_fft_64_stage_2_0_t409 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t946 = FSM_fft_64_stage_2_0_t945[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t947 = FSM_fft_64_stage_2_0_t946[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t948 = FSM_fft_64_stage_2_0_t927[FSM_fft_64_stage_2_0_t947 * 32 +: 32];
    FSM_fft_64_stage_2_0_t949 = FSM_fft_64_stage_2_0_t409 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t950 = FSM_fft_64_stage_2_0_t949[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t951 = FSM_fft_64_stage_2_0_t950[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t952 = FSM_fft_64_stage_2_0_t927[FSM_fft_64_stage_2_0_t951 * 32 +: 32];
    FSM_fft_64_stage_2_0_t953 = FSM_fft_64_stage_2_0_t948 + FSM_fft_64_stage_2_0_t952;
    FSM_fft_64_stage_2_0_t954 = FSM_fft_64_stage_2_0_t953[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t955 = FSM_fft_64_stage_2_0_t941;
    FSM_fft_64_stage_2_0_t955[FSM_fft_64_stage_2_0_t944 * 32 +: 32] = FSM_fft_64_stage_2_0_t954;
    FSM_fft_64_stage_2_0_t956 = FSM_fft_64_stage_2_0_t409 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t957 = FSM_fft_64_stage_2_0_t956[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t958 = FSM_fft_64_stage_2_0_t957[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t959 = FSM_fft_64_stage_2_0_t955;
    FSM_fft_64_stage_2_0_t959[FSM_fft_64_stage_2_0_t958 * 32 +: 32] = FSM_fft_64_stage_2_0_t948 - FSM_fft_64_stage_2_0_t952;
    FSM_fft_64_stage_2_0_t960 = FSM_fft_64_stage_2_0_t443[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t961 = FSM_fft_64_stage_2_0_t443[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t962 = FSM_fft_64_stage_2_0_t959[FSM_fft_64_stage_2_0_t961 * 32 +: 32];
    FSM_fft_64_stage_2_0_t963 = FSM_fft_64_stage_2_0_t443 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t964 = FSM_fft_64_stage_2_0_t963[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t965 = FSM_fft_64_stage_2_0_t964[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t966 = FSM_fft_64_stage_2_0_t959[FSM_fft_64_stage_2_0_t965 * 32 +: 32];
    FSM_fft_64_stage_2_0_t967 = FSM_fft_64_stage_2_0_t962 + FSM_fft_64_stage_2_0_t966;
    FSM_fft_64_stage_2_0_t968 = FSM_fft_64_stage_2_0_t967[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t969 = FSM_fft_64_stage_2_0_t959;
    FSM_fft_64_stage_2_0_t969[FSM_fft_64_stage_2_0_t960 * 32 +: 32] = FSM_fft_64_stage_2_0_t968;
    FSM_fft_64_stage_2_0_t970 = FSM_fft_64_stage_2_0_t443 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t971 = FSM_fft_64_stage_2_0_t970[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t972 = FSM_fft_64_stage_2_0_t971[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t973 = FSM_fft_64_stage_2_0_t969;
    FSM_fft_64_stage_2_0_t973[FSM_fft_64_stage_2_0_t972 * 32 +: 32] = FSM_fft_64_stage_2_0_t962 - FSM_fft_64_stage_2_0_t966;
    FSM_fft_64_stage_2_0_t974 = FSM_fft_64_stage_2_0_t443 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t975 = FSM_fft_64_stage_2_0_t974[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t976 = FSM_fft_64_stage_2_0_t975[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t977 = FSM_fft_64_stage_2_0_t443 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t978 = FSM_fft_64_stage_2_0_t977[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t979 = FSM_fft_64_stage_2_0_t978[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t980 = FSM_fft_64_stage_2_0_t959[FSM_fft_64_stage_2_0_t979 * 32 +: 32];
    FSM_fft_64_stage_2_0_t981 = FSM_fft_64_stage_2_0_t443 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t982 = FSM_fft_64_stage_2_0_t981[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t983 = FSM_fft_64_stage_2_0_t982[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t984 = FSM_fft_64_stage_2_0_t959[FSM_fft_64_stage_2_0_t983 * 32 +: 32];
    FSM_fft_64_stage_2_0_t985 = FSM_fft_64_stage_2_0_t980 + FSM_fft_64_stage_2_0_t984;
    FSM_fft_64_stage_2_0_t986 = FSM_fft_64_stage_2_0_t985[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t987 = FSM_fft_64_stage_2_0_t973;
    FSM_fft_64_stage_2_0_t987[FSM_fft_64_stage_2_0_t976 * 32 +: 32] = FSM_fft_64_stage_2_0_t986;
    FSM_fft_64_stage_2_0_t988 = FSM_fft_64_stage_2_0_t443 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t989 = FSM_fft_64_stage_2_0_t988[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t990 = FSM_fft_64_stage_2_0_t989[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t991 = FSM_fft_64_stage_2_0_t987;
    FSM_fft_64_stage_2_0_t991[FSM_fft_64_stage_2_0_t990 * 32 +: 32] = FSM_fft_64_stage_2_0_t980 - FSM_fft_64_stage_2_0_t984;
    FSM_fft_64_stage_2_0_t992 = FSM_fft_64_stage_2_0_t477[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t993 = FSM_fft_64_stage_2_0_t477[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t994 = FSM_fft_64_stage_2_0_t991[FSM_fft_64_stage_2_0_t993 * 32 +: 32];
    FSM_fft_64_stage_2_0_t995 = FSM_fft_64_stage_2_0_t477 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t996 = FSM_fft_64_stage_2_0_t995[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t997 = FSM_fft_64_stage_2_0_t996[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t998 = FSM_fft_64_stage_2_0_t991[FSM_fft_64_stage_2_0_t997 * 32 +: 32];
    FSM_fft_64_stage_2_0_t999 = FSM_fft_64_stage_2_0_t994 + FSM_fft_64_stage_2_0_t998;
    FSM_fft_64_stage_2_0_t1000 = FSM_fft_64_stage_2_0_t999[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t1001 = FSM_fft_64_stage_2_0_t991;
    FSM_fft_64_stage_2_0_t1001[FSM_fft_64_stage_2_0_t992 * 32 +: 32] = FSM_fft_64_stage_2_0_t1000;
    FSM_fft_64_stage_2_0_t1002 = FSM_fft_64_stage_2_0_t477 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t1003 = FSM_fft_64_stage_2_0_t1002[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t1004 = FSM_fft_64_stage_2_0_t1003[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t1005 = FSM_fft_64_stage_2_0_t1001;
    FSM_fft_64_stage_2_0_t1005[FSM_fft_64_stage_2_0_t1004 * 32 +: 32] = FSM_fft_64_stage_2_0_t994 - FSM_fft_64_stage_2_0_t998;
    FSM_fft_64_stage_2_0_t1006 = FSM_fft_64_stage_2_0_t477 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t1007 = FSM_fft_64_stage_2_0_t1006[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t1008 = FSM_fft_64_stage_2_0_t1007[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t1009 = FSM_fft_64_stage_2_0_t477 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t1010 = FSM_fft_64_stage_2_0_t1009[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t1011 = FSM_fft_64_stage_2_0_t1010[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t1012 = FSM_fft_64_stage_2_0_t991[FSM_fft_64_stage_2_0_t1011 * 32 +: 32];
    FSM_fft_64_stage_2_0_t1013 = FSM_fft_64_stage_2_0_t477 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t1014 = FSM_fft_64_stage_2_0_t1013[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t1015 = FSM_fft_64_stage_2_0_t1014[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t1016 = FSM_fft_64_stage_2_0_t991[FSM_fft_64_stage_2_0_t1015 * 32 +: 32];
    FSM_fft_64_stage_2_0_t1017 = FSM_fft_64_stage_2_0_t1012 + FSM_fft_64_stage_2_0_t1016;
    FSM_fft_64_stage_2_0_t1018 = FSM_fft_64_stage_2_0_t1017[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t1019 = FSM_fft_64_stage_2_0_t1005;
    FSM_fft_64_stage_2_0_t1019[FSM_fft_64_stage_2_0_t1008 * 32 +: 32] = FSM_fft_64_stage_2_0_t1018;
    FSM_fft_64_stage_2_0_t1020 = FSM_fft_64_stage_2_0_t477 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t1021 = FSM_fft_64_stage_2_0_t1020[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t1022 = FSM_fft_64_stage_2_0_t1021[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t1023 = FSM_fft_64_stage_2_0_t1019;
    FSM_fft_64_stage_2_0_t1023[FSM_fft_64_stage_2_0_t1022 * 32 +: 32] = FSM_fft_64_stage_2_0_t1012 - FSM_fft_64_stage_2_0_t1016;
    FSM_fft_64_stage_2_0_t1024 = FSM_fft_64_stage_2_0_t511[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t1025 = FSM_fft_64_stage_2_0_t511[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t1026 = FSM_fft_64_stage_2_0_t1023[FSM_fft_64_stage_2_0_t1025 * 32 +: 32];
    FSM_fft_64_stage_2_0_t1027 = FSM_fft_64_stage_2_0_t511 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t1028 = FSM_fft_64_stage_2_0_t1027[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t1029 = FSM_fft_64_stage_2_0_t1028[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t1030 = FSM_fft_64_stage_2_0_t1023[FSM_fft_64_stage_2_0_t1029 * 32 +: 32];
    FSM_fft_64_stage_2_0_t1031 = FSM_fft_64_stage_2_0_t1026 + FSM_fft_64_stage_2_0_t1030;
    FSM_fft_64_stage_2_0_t1032 = FSM_fft_64_stage_2_0_t1031[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t1033 = FSM_fft_64_stage_2_0_t1023;
    FSM_fft_64_stage_2_0_t1033[FSM_fft_64_stage_2_0_t1024 * 32 +: 32] = FSM_fft_64_stage_2_0_t1032;
    FSM_fft_64_stage_2_0_t1034 = FSM_fft_64_stage_2_0_t511 + 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_2_0_t1035 = FSM_fft_64_stage_2_0_t1034[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t1036 = FSM_fft_64_stage_2_0_t1035[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t1037 = FSM_fft_64_stage_2_0_t1033;
    FSM_fft_64_stage_2_0_t1037[FSM_fft_64_stage_2_0_t1036 * 32 +: 32] = FSM_fft_64_stage_2_0_t1026 - FSM_fft_64_stage_2_0_t1030;
    FSM_fft_64_stage_2_0_t1038 = FSM_fft_64_stage_2_0_t511 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t1039 = FSM_fft_64_stage_2_0_t1038[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t1040 = FSM_fft_64_stage_2_0_t1039[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t1041 = FSM_fft_64_stage_2_0_t511 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_2_0_t1042 = FSM_fft_64_stage_2_0_t1041[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t1043 = FSM_fft_64_stage_2_0_t1042[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t1044 = FSM_fft_64_stage_2_0_t1023[FSM_fft_64_stage_2_0_t1043 * 32 +: 32];
    FSM_fft_64_stage_2_0_t1045 = FSM_fft_64_stage_2_0_t511 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t1046 = FSM_fft_64_stage_2_0_t1045[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t1047 = FSM_fft_64_stage_2_0_t1046[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t1048 = FSM_fft_64_stage_2_0_t1023[FSM_fft_64_stage_2_0_t1047 * 32 +: 32];
    FSM_fft_64_stage_2_0_t1049 = FSM_fft_64_stage_2_0_t1044 + FSM_fft_64_stage_2_0_t1048;
    FSM_fft_64_stage_2_0_t1050 = FSM_fft_64_stage_2_0_t1049[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t1051 = FSM_fft_64_stage_2_0_t1037;
    FSM_fft_64_stage_2_0_t1051[FSM_fft_64_stage_2_0_t1040 * 32 +: 32] = FSM_fft_64_stage_2_0_t1050;
    FSM_fft_64_stage_2_0_t1052 = FSM_fft_64_stage_2_0_t511 + 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_2_0_t1053 = FSM_fft_64_stage_2_0_t1052[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_2_0_t1054 = FSM_fft_64_stage_2_0_t1053[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_2_0_t1055 = FSM_fft_64_stage_2_0_t1051;
    FSM_fft_64_stage_2_0_t1055[FSM_fft_64_stage_2_0_t1054 * 32 +: 32] = FSM_fft_64_stage_2_0_t1044 - FSM_fft_64_stage_2_0_t1048;
end

assign FSM_fft_64_stage_2_0_in_ready = 1'b1;

always @(posedge clk) begin
    FSM_fft_64_stage_2_0_st_dummy_reg <= FSM_fft_64_stage_2_0_st_dummy_reg;
    if (rst) begin
        FSM_fft_64_stage_2_0_st_dummy_reg <= 32'b0;
    end
end
/* End submodules of fft_64_stage_2 */
/* End module fft_64_stage_2 */
endgenerate
endmodule
