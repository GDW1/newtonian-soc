`timescale 1ns / 1ps

module fft_64_stage_1_inner
(
    input wire clk,
    input wire rst,
    input wire [2048-1:0] i_data_in_real,
    input wire [2048-1:0] i_data_in_imag,
    input wire i_valid,
    output wire i_ready,
    output wire [2048-1:0] o_data_out_real,
    output wire [2048-1:0] o_data_out_imag,
    output wire o_valid,
    input wire o_ready
);

generate
/*
    Begin module fft_64_stage_1
*/
/*
    Wires declared by fft_64_stage_1
*/
wire FSM_fft_64_stage_1_0_in_ready;
wire FSM_fft_64_stage_1_0_out_valid;
/* End wires declared by fft_64_stage_1 */

/*
    Submodules of fft_64_stage_1
*/
reg [32-1:0] FSM_fft_64_stage_1_0_st_dummy_reg = 32'b0;

reg [64-1:0] FSM_fft_64_stage_1_0_t0;
reg [32-1:0] FSM_fft_64_stage_1_0_t1;
reg [6-1:0] FSM_fft_64_stage_1_0_t2;
reg [64-1:0] FSM_fft_64_stage_1_0_t3;
reg [32-1:0] FSM_fft_64_stage_1_0_t4;
reg [6-1:0] FSM_fft_64_stage_1_0_t5;
reg [32-1:0] FSM_fft_64_stage_1_0_t6;
reg [64-1:0] FSM_fft_64_stage_1_0_t7;
reg [32-1:0] FSM_fft_64_stage_1_0_t8;
reg [33-1:0] FSM_fft_64_stage_1_0_t9;
reg [32-1:0] FSM_fft_64_stage_1_0_t10;
reg [6-1:0] FSM_fft_64_stage_1_0_t11;
reg [32-1:0] FSM_fft_64_stage_1_0_t12;
reg [33-1:0] FSM_fft_64_stage_1_0_t13;
reg [32-1:0] FSM_fft_64_stage_1_0_t14;
reg [2048-1:0] FSM_fft_64_stage_1_0_t15;
reg [64-1:0] FSM_fft_64_stage_1_0_t16;
reg [32-1:0] FSM_fft_64_stage_1_0_t17;
reg [33-1:0] FSM_fft_64_stage_1_0_t18;
reg [32-1:0] FSM_fft_64_stage_1_0_t19;
reg [6-1:0] FSM_fft_64_stage_1_0_t20;
reg [2048-1:0] FSM_fft_64_stage_1_0_t21;
reg [64-1:0] FSM_fft_64_stage_1_0_t22;
reg [32-1:0] FSM_fft_64_stage_1_0_t23;
reg [6-1:0] FSM_fft_64_stage_1_0_t24;
reg [64-1:0] FSM_fft_64_stage_1_0_t25;
reg [32-1:0] FSM_fft_64_stage_1_0_t26;
reg [6-1:0] FSM_fft_64_stage_1_0_t27;
reg [32-1:0] FSM_fft_64_stage_1_0_t28;
reg [64-1:0] FSM_fft_64_stage_1_0_t29;
reg [32-1:0] FSM_fft_64_stage_1_0_t30;
reg [33-1:0] FSM_fft_64_stage_1_0_t31;
reg [32-1:0] FSM_fft_64_stage_1_0_t32;
reg [6-1:0] FSM_fft_64_stage_1_0_t33;
reg [32-1:0] FSM_fft_64_stage_1_0_t34;
reg [33-1:0] FSM_fft_64_stage_1_0_t35;
reg [32-1:0] FSM_fft_64_stage_1_0_t36;
reg [2048-1:0] FSM_fft_64_stage_1_0_t37;
reg [64-1:0] FSM_fft_64_stage_1_0_t38;
reg [32-1:0] FSM_fft_64_stage_1_0_t39;
reg [33-1:0] FSM_fft_64_stage_1_0_t40;
reg [32-1:0] FSM_fft_64_stage_1_0_t41;
reg [6-1:0] FSM_fft_64_stage_1_0_t42;
reg [2048-1:0] FSM_fft_64_stage_1_0_t43;
reg [64-1:0] FSM_fft_64_stage_1_0_t44;
reg [32-1:0] FSM_fft_64_stage_1_0_t45;
reg [6-1:0] FSM_fft_64_stage_1_0_t46;
reg [64-1:0] FSM_fft_64_stage_1_0_t47;
reg [32-1:0] FSM_fft_64_stage_1_0_t48;
reg [6-1:0] FSM_fft_64_stage_1_0_t49;
reg [32-1:0] FSM_fft_64_stage_1_0_t50;
reg [64-1:0] FSM_fft_64_stage_1_0_t51;
reg [32-1:0] FSM_fft_64_stage_1_0_t52;
reg [33-1:0] FSM_fft_64_stage_1_0_t53;
reg [32-1:0] FSM_fft_64_stage_1_0_t54;
reg [6-1:0] FSM_fft_64_stage_1_0_t55;
reg [32-1:0] FSM_fft_64_stage_1_0_t56;
reg [33-1:0] FSM_fft_64_stage_1_0_t57;
reg [32-1:0] FSM_fft_64_stage_1_0_t58;
reg [2048-1:0] FSM_fft_64_stage_1_0_t59;
reg [64-1:0] FSM_fft_64_stage_1_0_t60;
reg [32-1:0] FSM_fft_64_stage_1_0_t61;
reg [33-1:0] FSM_fft_64_stage_1_0_t62;
reg [32-1:0] FSM_fft_64_stage_1_0_t63;
reg [6-1:0] FSM_fft_64_stage_1_0_t64;
reg [2048-1:0] FSM_fft_64_stage_1_0_t65;
reg [64-1:0] FSM_fft_64_stage_1_0_t66;
reg [32-1:0] FSM_fft_64_stage_1_0_t67;
reg [6-1:0] FSM_fft_64_stage_1_0_t68;
reg [64-1:0] FSM_fft_64_stage_1_0_t69;
reg [32-1:0] FSM_fft_64_stage_1_0_t70;
reg [6-1:0] FSM_fft_64_stage_1_0_t71;
reg [32-1:0] FSM_fft_64_stage_1_0_t72;
reg [64-1:0] FSM_fft_64_stage_1_0_t73;
reg [32-1:0] FSM_fft_64_stage_1_0_t74;
reg [33-1:0] FSM_fft_64_stage_1_0_t75;
reg [32-1:0] FSM_fft_64_stage_1_0_t76;
reg [6-1:0] FSM_fft_64_stage_1_0_t77;
reg [32-1:0] FSM_fft_64_stage_1_0_t78;
reg [33-1:0] FSM_fft_64_stage_1_0_t79;
reg [32-1:0] FSM_fft_64_stage_1_0_t80;
reg [2048-1:0] FSM_fft_64_stage_1_0_t81;
reg [64-1:0] FSM_fft_64_stage_1_0_t82;
reg [32-1:0] FSM_fft_64_stage_1_0_t83;
reg [33-1:0] FSM_fft_64_stage_1_0_t84;
reg [32-1:0] FSM_fft_64_stage_1_0_t85;
reg [6-1:0] FSM_fft_64_stage_1_0_t86;
reg [2048-1:0] FSM_fft_64_stage_1_0_t87;
reg [64-1:0] FSM_fft_64_stage_1_0_t88;
reg [32-1:0] FSM_fft_64_stage_1_0_t89;
reg [6-1:0] FSM_fft_64_stage_1_0_t90;
reg [64-1:0] FSM_fft_64_stage_1_0_t91;
reg [32-1:0] FSM_fft_64_stage_1_0_t92;
reg [6-1:0] FSM_fft_64_stage_1_0_t93;
reg [32-1:0] FSM_fft_64_stage_1_0_t94;
reg [64-1:0] FSM_fft_64_stage_1_0_t95;
reg [32-1:0] FSM_fft_64_stage_1_0_t96;
reg [33-1:0] FSM_fft_64_stage_1_0_t97;
reg [32-1:0] FSM_fft_64_stage_1_0_t98;
reg [6-1:0] FSM_fft_64_stage_1_0_t99;
reg [32-1:0] FSM_fft_64_stage_1_0_t100;
reg [33-1:0] FSM_fft_64_stage_1_0_t101;
reg [32-1:0] FSM_fft_64_stage_1_0_t102;
reg [2048-1:0] FSM_fft_64_stage_1_0_t103;
reg [64-1:0] FSM_fft_64_stage_1_0_t104;
reg [32-1:0] FSM_fft_64_stage_1_0_t105;
reg [33-1:0] FSM_fft_64_stage_1_0_t106;
reg [32-1:0] FSM_fft_64_stage_1_0_t107;
reg [6-1:0] FSM_fft_64_stage_1_0_t108;
reg [2048-1:0] FSM_fft_64_stage_1_0_t109;
reg [64-1:0] FSM_fft_64_stage_1_0_t110;
reg [32-1:0] FSM_fft_64_stage_1_0_t111;
reg [6-1:0] FSM_fft_64_stage_1_0_t112;
reg [64-1:0] FSM_fft_64_stage_1_0_t113;
reg [32-1:0] FSM_fft_64_stage_1_0_t114;
reg [6-1:0] FSM_fft_64_stage_1_0_t115;
reg [32-1:0] FSM_fft_64_stage_1_0_t116;
reg [64-1:0] FSM_fft_64_stage_1_0_t117;
reg [32-1:0] FSM_fft_64_stage_1_0_t118;
reg [33-1:0] FSM_fft_64_stage_1_0_t119;
reg [32-1:0] FSM_fft_64_stage_1_0_t120;
reg [6-1:0] FSM_fft_64_stage_1_0_t121;
reg [32-1:0] FSM_fft_64_stage_1_0_t122;
reg [33-1:0] FSM_fft_64_stage_1_0_t123;
reg [32-1:0] FSM_fft_64_stage_1_0_t124;
reg [2048-1:0] FSM_fft_64_stage_1_0_t125;
reg [64-1:0] FSM_fft_64_stage_1_0_t126;
reg [32-1:0] FSM_fft_64_stage_1_0_t127;
reg [33-1:0] FSM_fft_64_stage_1_0_t128;
reg [32-1:0] FSM_fft_64_stage_1_0_t129;
reg [6-1:0] FSM_fft_64_stage_1_0_t130;
reg [2048-1:0] FSM_fft_64_stage_1_0_t131;
reg [64-1:0] FSM_fft_64_stage_1_0_t132;
reg [32-1:0] FSM_fft_64_stage_1_0_t133;
reg [6-1:0] FSM_fft_64_stage_1_0_t134;
reg [64-1:0] FSM_fft_64_stage_1_0_t135;
reg [32-1:0] FSM_fft_64_stage_1_0_t136;
reg [6-1:0] FSM_fft_64_stage_1_0_t137;
reg [32-1:0] FSM_fft_64_stage_1_0_t138;
reg [64-1:0] FSM_fft_64_stage_1_0_t139;
reg [32-1:0] FSM_fft_64_stage_1_0_t140;
reg [33-1:0] FSM_fft_64_stage_1_0_t141;
reg [32-1:0] FSM_fft_64_stage_1_0_t142;
reg [6-1:0] FSM_fft_64_stage_1_0_t143;
reg [32-1:0] FSM_fft_64_stage_1_0_t144;
reg [33-1:0] FSM_fft_64_stage_1_0_t145;
reg [32-1:0] FSM_fft_64_stage_1_0_t146;
reg [2048-1:0] FSM_fft_64_stage_1_0_t147;
reg [64-1:0] FSM_fft_64_stage_1_0_t148;
reg [32-1:0] FSM_fft_64_stage_1_0_t149;
reg [33-1:0] FSM_fft_64_stage_1_0_t150;
reg [32-1:0] FSM_fft_64_stage_1_0_t151;
reg [6-1:0] FSM_fft_64_stage_1_0_t152;
reg [2048-1:0] FSM_fft_64_stage_1_0_t153;
reg [64-1:0] FSM_fft_64_stage_1_0_t154;
reg [32-1:0] FSM_fft_64_stage_1_0_t155;
reg [6-1:0] FSM_fft_64_stage_1_0_t156;
reg [64-1:0] FSM_fft_64_stage_1_0_t157;
reg [32-1:0] FSM_fft_64_stage_1_0_t158;
reg [6-1:0] FSM_fft_64_stage_1_0_t159;
reg [32-1:0] FSM_fft_64_stage_1_0_t160;
reg [64-1:0] FSM_fft_64_stage_1_0_t161;
reg [32-1:0] FSM_fft_64_stage_1_0_t162;
reg [33-1:0] FSM_fft_64_stage_1_0_t163;
reg [32-1:0] FSM_fft_64_stage_1_0_t164;
reg [6-1:0] FSM_fft_64_stage_1_0_t165;
reg [32-1:0] FSM_fft_64_stage_1_0_t166;
reg [33-1:0] FSM_fft_64_stage_1_0_t167;
reg [32-1:0] FSM_fft_64_stage_1_0_t168;
reg [2048-1:0] FSM_fft_64_stage_1_0_t169;
reg [64-1:0] FSM_fft_64_stage_1_0_t170;
reg [32-1:0] FSM_fft_64_stage_1_0_t171;
reg [33-1:0] FSM_fft_64_stage_1_0_t172;
reg [32-1:0] FSM_fft_64_stage_1_0_t173;
reg [6-1:0] FSM_fft_64_stage_1_0_t174;
reg [2048-1:0] FSM_fft_64_stage_1_0_t175;
reg [64-1:0] FSM_fft_64_stage_1_0_t176;
reg [32-1:0] FSM_fft_64_stage_1_0_t177;
reg [6-1:0] FSM_fft_64_stage_1_0_t178;
reg [64-1:0] FSM_fft_64_stage_1_0_t179;
reg [32-1:0] FSM_fft_64_stage_1_0_t180;
reg [6-1:0] FSM_fft_64_stage_1_0_t181;
reg [32-1:0] FSM_fft_64_stage_1_0_t182;
reg [64-1:0] FSM_fft_64_stage_1_0_t183;
reg [32-1:0] FSM_fft_64_stage_1_0_t184;
reg [33-1:0] FSM_fft_64_stage_1_0_t185;
reg [32-1:0] FSM_fft_64_stage_1_0_t186;
reg [6-1:0] FSM_fft_64_stage_1_0_t187;
reg [32-1:0] FSM_fft_64_stage_1_0_t188;
reg [33-1:0] FSM_fft_64_stage_1_0_t189;
reg [32-1:0] FSM_fft_64_stage_1_0_t190;
reg [2048-1:0] FSM_fft_64_stage_1_0_t191;
reg [64-1:0] FSM_fft_64_stage_1_0_t192;
reg [32-1:0] FSM_fft_64_stage_1_0_t193;
reg [33-1:0] FSM_fft_64_stage_1_0_t194;
reg [32-1:0] FSM_fft_64_stage_1_0_t195;
reg [6-1:0] FSM_fft_64_stage_1_0_t196;
reg [2048-1:0] FSM_fft_64_stage_1_0_t197;
reg [64-1:0] FSM_fft_64_stage_1_0_t198;
reg [32-1:0] FSM_fft_64_stage_1_0_t199;
reg [6-1:0] FSM_fft_64_stage_1_0_t200;
reg [64-1:0] FSM_fft_64_stage_1_0_t201;
reg [32-1:0] FSM_fft_64_stage_1_0_t202;
reg [6-1:0] FSM_fft_64_stage_1_0_t203;
reg [32-1:0] FSM_fft_64_stage_1_0_t204;
reg [64-1:0] FSM_fft_64_stage_1_0_t205;
reg [32-1:0] FSM_fft_64_stage_1_0_t206;
reg [33-1:0] FSM_fft_64_stage_1_0_t207;
reg [32-1:0] FSM_fft_64_stage_1_0_t208;
reg [6-1:0] FSM_fft_64_stage_1_0_t209;
reg [32-1:0] FSM_fft_64_stage_1_0_t210;
reg [33-1:0] FSM_fft_64_stage_1_0_t211;
reg [32-1:0] FSM_fft_64_stage_1_0_t212;
reg [2048-1:0] FSM_fft_64_stage_1_0_t213;
reg [64-1:0] FSM_fft_64_stage_1_0_t214;
reg [32-1:0] FSM_fft_64_stage_1_0_t215;
reg [33-1:0] FSM_fft_64_stage_1_0_t216;
reg [32-1:0] FSM_fft_64_stage_1_0_t217;
reg [6-1:0] FSM_fft_64_stage_1_0_t218;
reg [2048-1:0] FSM_fft_64_stage_1_0_t219;
reg [64-1:0] FSM_fft_64_stage_1_0_t220;
reg [32-1:0] FSM_fft_64_stage_1_0_t221;
reg [6-1:0] FSM_fft_64_stage_1_0_t222;
reg [64-1:0] FSM_fft_64_stage_1_0_t223;
reg [32-1:0] FSM_fft_64_stage_1_0_t224;
reg [6-1:0] FSM_fft_64_stage_1_0_t225;
reg [32-1:0] FSM_fft_64_stage_1_0_t226;
reg [64-1:0] FSM_fft_64_stage_1_0_t227;
reg [32-1:0] FSM_fft_64_stage_1_0_t228;
reg [33-1:0] FSM_fft_64_stage_1_0_t229;
reg [32-1:0] FSM_fft_64_stage_1_0_t230;
reg [6-1:0] FSM_fft_64_stage_1_0_t231;
reg [32-1:0] FSM_fft_64_stage_1_0_t232;
reg [33-1:0] FSM_fft_64_stage_1_0_t233;
reg [32-1:0] FSM_fft_64_stage_1_0_t234;
reg [2048-1:0] FSM_fft_64_stage_1_0_t235;
reg [64-1:0] FSM_fft_64_stage_1_0_t236;
reg [32-1:0] FSM_fft_64_stage_1_0_t237;
reg [33-1:0] FSM_fft_64_stage_1_0_t238;
reg [32-1:0] FSM_fft_64_stage_1_0_t239;
reg [6-1:0] FSM_fft_64_stage_1_0_t240;
reg [2048-1:0] FSM_fft_64_stage_1_0_t241;
reg [64-1:0] FSM_fft_64_stage_1_0_t242;
reg [32-1:0] FSM_fft_64_stage_1_0_t243;
reg [6-1:0] FSM_fft_64_stage_1_0_t244;
reg [64-1:0] FSM_fft_64_stage_1_0_t245;
reg [32-1:0] FSM_fft_64_stage_1_0_t246;
reg [6-1:0] FSM_fft_64_stage_1_0_t247;
reg [32-1:0] FSM_fft_64_stage_1_0_t248;
reg [64-1:0] FSM_fft_64_stage_1_0_t249;
reg [32-1:0] FSM_fft_64_stage_1_0_t250;
reg [33-1:0] FSM_fft_64_stage_1_0_t251;
reg [32-1:0] FSM_fft_64_stage_1_0_t252;
reg [6-1:0] FSM_fft_64_stage_1_0_t253;
reg [32-1:0] FSM_fft_64_stage_1_0_t254;
reg [33-1:0] FSM_fft_64_stage_1_0_t255;
reg [32-1:0] FSM_fft_64_stage_1_0_t256;
reg [2048-1:0] FSM_fft_64_stage_1_0_t257;
reg [64-1:0] FSM_fft_64_stage_1_0_t258;
reg [32-1:0] FSM_fft_64_stage_1_0_t259;
reg [33-1:0] FSM_fft_64_stage_1_0_t260;
reg [32-1:0] FSM_fft_64_stage_1_0_t261;
reg [6-1:0] FSM_fft_64_stage_1_0_t262;
reg [2048-1:0] FSM_fft_64_stage_1_0_t263;
reg [64-1:0] FSM_fft_64_stage_1_0_t264;
reg [32-1:0] FSM_fft_64_stage_1_0_t265;
reg [6-1:0] FSM_fft_64_stage_1_0_t266;
reg [64-1:0] FSM_fft_64_stage_1_0_t267;
reg [32-1:0] FSM_fft_64_stage_1_0_t268;
reg [6-1:0] FSM_fft_64_stage_1_0_t269;
reg [32-1:0] FSM_fft_64_stage_1_0_t270;
reg [64-1:0] FSM_fft_64_stage_1_0_t271;
reg [32-1:0] FSM_fft_64_stage_1_0_t272;
reg [33-1:0] FSM_fft_64_stage_1_0_t273;
reg [32-1:0] FSM_fft_64_stage_1_0_t274;
reg [6-1:0] FSM_fft_64_stage_1_0_t275;
reg [32-1:0] FSM_fft_64_stage_1_0_t276;
reg [33-1:0] FSM_fft_64_stage_1_0_t277;
reg [32-1:0] FSM_fft_64_stage_1_0_t278;
reg [2048-1:0] FSM_fft_64_stage_1_0_t279;
reg [64-1:0] FSM_fft_64_stage_1_0_t280;
reg [32-1:0] FSM_fft_64_stage_1_0_t281;
reg [33-1:0] FSM_fft_64_stage_1_0_t282;
reg [32-1:0] FSM_fft_64_stage_1_0_t283;
reg [6-1:0] FSM_fft_64_stage_1_0_t284;
reg [2048-1:0] FSM_fft_64_stage_1_0_t285;
reg [64-1:0] FSM_fft_64_stage_1_0_t286;
reg [32-1:0] FSM_fft_64_stage_1_0_t287;
reg [6-1:0] FSM_fft_64_stage_1_0_t288;
reg [64-1:0] FSM_fft_64_stage_1_0_t289;
reg [32-1:0] FSM_fft_64_stage_1_0_t290;
reg [6-1:0] FSM_fft_64_stage_1_0_t291;
reg [32-1:0] FSM_fft_64_stage_1_0_t292;
reg [64-1:0] FSM_fft_64_stage_1_0_t293;
reg [32-1:0] FSM_fft_64_stage_1_0_t294;
reg [33-1:0] FSM_fft_64_stage_1_0_t295;
reg [32-1:0] FSM_fft_64_stage_1_0_t296;
reg [6-1:0] FSM_fft_64_stage_1_0_t297;
reg [32-1:0] FSM_fft_64_stage_1_0_t298;
reg [33-1:0] FSM_fft_64_stage_1_0_t299;
reg [32-1:0] FSM_fft_64_stage_1_0_t300;
reg [2048-1:0] FSM_fft_64_stage_1_0_t301;
reg [64-1:0] FSM_fft_64_stage_1_0_t302;
reg [32-1:0] FSM_fft_64_stage_1_0_t303;
reg [33-1:0] FSM_fft_64_stage_1_0_t304;
reg [32-1:0] FSM_fft_64_stage_1_0_t305;
reg [6-1:0] FSM_fft_64_stage_1_0_t306;
reg [2048-1:0] FSM_fft_64_stage_1_0_t307;
reg [64-1:0] FSM_fft_64_stage_1_0_t308;
reg [32-1:0] FSM_fft_64_stage_1_0_t309;
reg [6-1:0] FSM_fft_64_stage_1_0_t310;
reg [64-1:0] FSM_fft_64_stage_1_0_t311;
reg [32-1:0] FSM_fft_64_stage_1_0_t312;
reg [6-1:0] FSM_fft_64_stage_1_0_t313;
reg [32-1:0] FSM_fft_64_stage_1_0_t314;
reg [64-1:0] FSM_fft_64_stage_1_0_t315;
reg [32-1:0] FSM_fft_64_stage_1_0_t316;
reg [33-1:0] FSM_fft_64_stage_1_0_t317;
reg [32-1:0] FSM_fft_64_stage_1_0_t318;
reg [6-1:0] FSM_fft_64_stage_1_0_t319;
reg [32-1:0] FSM_fft_64_stage_1_0_t320;
reg [33-1:0] FSM_fft_64_stage_1_0_t321;
reg [32-1:0] FSM_fft_64_stage_1_0_t322;
reg [2048-1:0] FSM_fft_64_stage_1_0_t323;
reg [64-1:0] FSM_fft_64_stage_1_0_t324;
reg [32-1:0] FSM_fft_64_stage_1_0_t325;
reg [33-1:0] FSM_fft_64_stage_1_0_t326;
reg [32-1:0] FSM_fft_64_stage_1_0_t327;
reg [6-1:0] FSM_fft_64_stage_1_0_t328;
reg [2048-1:0] FSM_fft_64_stage_1_0_t329;
reg [64-1:0] FSM_fft_64_stage_1_0_t330;
reg [32-1:0] FSM_fft_64_stage_1_0_t331;
reg [6-1:0] FSM_fft_64_stage_1_0_t332;
reg [64-1:0] FSM_fft_64_stage_1_0_t333;
reg [32-1:0] FSM_fft_64_stage_1_0_t334;
reg [6-1:0] FSM_fft_64_stage_1_0_t335;
reg [32-1:0] FSM_fft_64_stage_1_0_t336;
reg [64-1:0] FSM_fft_64_stage_1_0_t337;
reg [32-1:0] FSM_fft_64_stage_1_0_t338;
reg [33-1:0] FSM_fft_64_stage_1_0_t339;
reg [32-1:0] FSM_fft_64_stage_1_0_t340;
reg [6-1:0] FSM_fft_64_stage_1_0_t341;
reg [32-1:0] FSM_fft_64_stage_1_0_t342;
reg [33-1:0] FSM_fft_64_stage_1_0_t343;
reg [32-1:0] FSM_fft_64_stage_1_0_t344;
reg [2048-1:0] FSM_fft_64_stage_1_0_t345;
reg [64-1:0] FSM_fft_64_stage_1_0_t346;
reg [32-1:0] FSM_fft_64_stage_1_0_t347;
reg [33-1:0] FSM_fft_64_stage_1_0_t348;
reg [32-1:0] FSM_fft_64_stage_1_0_t349;
reg [6-1:0] FSM_fft_64_stage_1_0_t350;
reg [2048-1:0] FSM_fft_64_stage_1_0_t351;
reg [64-1:0] FSM_fft_64_stage_1_0_t352;
reg [32-1:0] FSM_fft_64_stage_1_0_t353;
reg [6-1:0] FSM_fft_64_stage_1_0_t354;
reg [64-1:0] FSM_fft_64_stage_1_0_t355;
reg [32-1:0] FSM_fft_64_stage_1_0_t356;
reg [6-1:0] FSM_fft_64_stage_1_0_t357;
reg [32-1:0] FSM_fft_64_stage_1_0_t358;
reg [64-1:0] FSM_fft_64_stage_1_0_t359;
reg [32-1:0] FSM_fft_64_stage_1_0_t360;
reg [33-1:0] FSM_fft_64_stage_1_0_t361;
reg [32-1:0] FSM_fft_64_stage_1_0_t362;
reg [6-1:0] FSM_fft_64_stage_1_0_t363;
reg [32-1:0] FSM_fft_64_stage_1_0_t364;
reg [33-1:0] FSM_fft_64_stage_1_0_t365;
reg [32-1:0] FSM_fft_64_stage_1_0_t366;
reg [2048-1:0] FSM_fft_64_stage_1_0_t367;
reg [64-1:0] FSM_fft_64_stage_1_0_t368;
reg [32-1:0] FSM_fft_64_stage_1_0_t369;
reg [33-1:0] FSM_fft_64_stage_1_0_t370;
reg [32-1:0] FSM_fft_64_stage_1_0_t371;
reg [6-1:0] FSM_fft_64_stage_1_0_t372;
reg [2048-1:0] FSM_fft_64_stage_1_0_t373;
reg [64-1:0] FSM_fft_64_stage_1_0_t374;
reg [32-1:0] FSM_fft_64_stage_1_0_t375;
reg [6-1:0] FSM_fft_64_stage_1_0_t376;
reg [64-1:0] FSM_fft_64_stage_1_0_t377;
reg [32-1:0] FSM_fft_64_stage_1_0_t378;
reg [6-1:0] FSM_fft_64_stage_1_0_t379;
reg [32-1:0] FSM_fft_64_stage_1_0_t380;
reg [64-1:0] FSM_fft_64_stage_1_0_t381;
reg [32-1:0] FSM_fft_64_stage_1_0_t382;
reg [33-1:0] FSM_fft_64_stage_1_0_t383;
reg [32-1:0] FSM_fft_64_stage_1_0_t384;
reg [6-1:0] FSM_fft_64_stage_1_0_t385;
reg [32-1:0] FSM_fft_64_stage_1_0_t386;
reg [33-1:0] FSM_fft_64_stage_1_0_t387;
reg [32-1:0] FSM_fft_64_stage_1_0_t388;
reg [2048-1:0] FSM_fft_64_stage_1_0_t389;
reg [64-1:0] FSM_fft_64_stage_1_0_t390;
reg [32-1:0] FSM_fft_64_stage_1_0_t391;
reg [33-1:0] FSM_fft_64_stage_1_0_t392;
reg [32-1:0] FSM_fft_64_stage_1_0_t393;
reg [6-1:0] FSM_fft_64_stage_1_0_t394;
reg [2048-1:0] FSM_fft_64_stage_1_0_t395;
reg [64-1:0] FSM_fft_64_stage_1_0_t396;
reg [32-1:0] FSM_fft_64_stage_1_0_t397;
reg [6-1:0] FSM_fft_64_stage_1_0_t398;
reg [64-1:0] FSM_fft_64_stage_1_0_t399;
reg [32-1:0] FSM_fft_64_stage_1_0_t400;
reg [6-1:0] FSM_fft_64_stage_1_0_t401;
reg [32-1:0] FSM_fft_64_stage_1_0_t402;
reg [64-1:0] FSM_fft_64_stage_1_0_t403;
reg [32-1:0] FSM_fft_64_stage_1_0_t404;
reg [33-1:0] FSM_fft_64_stage_1_0_t405;
reg [32-1:0] FSM_fft_64_stage_1_0_t406;
reg [6-1:0] FSM_fft_64_stage_1_0_t407;
reg [32-1:0] FSM_fft_64_stage_1_0_t408;
reg [33-1:0] FSM_fft_64_stage_1_0_t409;
reg [32-1:0] FSM_fft_64_stage_1_0_t410;
reg [2048-1:0] FSM_fft_64_stage_1_0_t411;
reg [64-1:0] FSM_fft_64_stage_1_0_t412;
reg [32-1:0] FSM_fft_64_stage_1_0_t413;
reg [33-1:0] FSM_fft_64_stage_1_0_t414;
reg [32-1:0] FSM_fft_64_stage_1_0_t415;
reg [6-1:0] FSM_fft_64_stage_1_0_t416;
reg [2048-1:0] FSM_fft_64_stage_1_0_t417;
reg [64-1:0] FSM_fft_64_stage_1_0_t418;
reg [32-1:0] FSM_fft_64_stage_1_0_t419;
reg [6-1:0] FSM_fft_64_stage_1_0_t420;
reg [64-1:0] FSM_fft_64_stage_1_0_t421;
reg [32-1:0] FSM_fft_64_stage_1_0_t422;
reg [6-1:0] FSM_fft_64_stage_1_0_t423;
reg [32-1:0] FSM_fft_64_stage_1_0_t424;
reg [64-1:0] FSM_fft_64_stage_1_0_t425;
reg [32-1:0] FSM_fft_64_stage_1_0_t426;
reg [33-1:0] FSM_fft_64_stage_1_0_t427;
reg [32-1:0] FSM_fft_64_stage_1_0_t428;
reg [6-1:0] FSM_fft_64_stage_1_0_t429;
reg [32-1:0] FSM_fft_64_stage_1_0_t430;
reg [33-1:0] FSM_fft_64_stage_1_0_t431;
reg [32-1:0] FSM_fft_64_stage_1_0_t432;
reg [2048-1:0] FSM_fft_64_stage_1_0_t433;
reg [64-1:0] FSM_fft_64_stage_1_0_t434;
reg [32-1:0] FSM_fft_64_stage_1_0_t435;
reg [33-1:0] FSM_fft_64_stage_1_0_t436;
reg [32-1:0] FSM_fft_64_stage_1_0_t437;
reg [6-1:0] FSM_fft_64_stage_1_0_t438;
reg [2048-1:0] FSM_fft_64_stage_1_0_t439;
reg [64-1:0] FSM_fft_64_stage_1_0_t440;
reg [32-1:0] FSM_fft_64_stage_1_0_t441;
reg [6-1:0] FSM_fft_64_stage_1_0_t442;
reg [64-1:0] FSM_fft_64_stage_1_0_t443;
reg [32-1:0] FSM_fft_64_stage_1_0_t444;
reg [6-1:0] FSM_fft_64_stage_1_0_t445;
reg [32-1:0] FSM_fft_64_stage_1_0_t446;
reg [64-1:0] FSM_fft_64_stage_1_0_t447;
reg [32-1:0] FSM_fft_64_stage_1_0_t448;
reg [33-1:0] FSM_fft_64_stage_1_0_t449;
reg [32-1:0] FSM_fft_64_stage_1_0_t450;
reg [6-1:0] FSM_fft_64_stage_1_0_t451;
reg [32-1:0] FSM_fft_64_stage_1_0_t452;
reg [33-1:0] FSM_fft_64_stage_1_0_t453;
reg [32-1:0] FSM_fft_64_stage_1_0_t454;
reg [2048-1:0] FSM_fft_64_stage_1_0_t455;
reg [64-1:0] FSM_fft_64_stage_1_0_t456;
reg [32-1:0] FSM_fft_64_stage_1_0_t457;
reg [33-1:0] FSM_fft_64_stage_1_0_t458;
reg [32-1:0] FSM_fft_64_stage_1_0_t459;
reg [6-1:0] FSM_fft_64_stage_1_0_t460;
reg [2048-1:0] FSM_fft_64_stage_1_0_t461;
reg [64-1:0] FSM_fft_64_stage_1_0_t462;
reg [32-1:0] FSM_fft_64_stage_1_0_t463;
reg [6-1:0] FSM_fft_64_stage_1_0_t464;
reg [64-1:0] FSM_fft_64_stage_1_0_t465;
reg [32-1:0] FSM_fft_64_stage_1_0_t466;
reg [6-1:0] FSM_fft_64_stage_1_0_t467;
reg [32-1:0] FSM_fft_64_stage_1_0_t468;
reg [64-1:0] FSM_fft_64_stage_1_0_t469;
reg [32-1:0] FSM_fft_64_stage_1_0_t470;
reg [33-1:0] FSM_fft_64_stage_1_0_t471;
reg [32-1:0] FSM_fft_64_stage_1_0_t472;
reg [6-1:0] FSM_fft_64_stage_1_0_t473;
reg [32-1:0] FSM_fft_64_stage_1_0_t474;
reg [33-1:0] FSM_fft_64_stage_1_0_t475;
reg [32-1:0] FSM_fft_64_stage_1_0_t476;
reg [2048-1:0] FSM_fft_64_stage_1_0_t477;
reg [64-1:0] FSM_fft_64_stage_1_0_t478;
reg [32-1:0] FSM_fft_64_stage_1_0_t479;
reg [33-1:0] FSM_fft_64_stage_1_0_t480;
reg [32-1:0] FSM_fft_64_stage_1_0_t481;
reg [6-1:0] FSM_fft_64_stage_1_0_t482;
reg [2048-1:0] FSM_fft_64_stage_1_0_t483;
reg [64-1:0] FSM_fft_64_stage_1_0_t484;
reg [32-1:0] FSM_fft_64_stage_1_0_t485;
reg [6-1:0] FSM_fft_64_stage_1_0_t486;
reg [64-1:0] FSM_fft_64_stage_1_0_t487;
reg [32-1:0] FSM_fft_64_stage_1_0_t488;
reg [6-1:0] FSM_fft_64_stage_1_0_t489;
reg [32-1:0] FSM_fft_64_stage_1_0_t490;
reg [64-1:0] FSM_fft_64_stage_1_0_t491;
reg [32-1:0] FSM_fft_64_stage_1_0_t492;
reg [33-1:0] FSM_fft_64_stage_1_0_t493;
reg [32-1:0] FSM_fft_64_stage_1_0_t494;
reg [6-1:0] FSM_fft_64_stage_1_0_t495;
reg [32-1:0] FSM_fft_64_stage_1_0_t496;
reg [33-1:0] FSM_fft_64_stage_1_0_t497;
reg [32-1:0] FSM_fft_64_stage_1_0_t498;
reg [2048-1:0] FSM_fft_64_stage_1_0_t499;
reg [64-1:0] FSM_fft_64_stage_1_0_t500;
reg [32-1:0] FSM_fft_64_stage_1_0_t501;
reg [33-1:0] FSM_fft_64_stage_1_0_t502;
reg [32-1:0] FSM_fft_64_stage_1_0_t503;
reg [6-1:0] FSM_fft_64_stage_1_0_t504;
reg [2048-1:0] FSM_fft_64_stage_1_0_t505;
reg [64-1:0] FSM_fft_64_stage_1_0_t506;
reg [32-1:0] FSM_fft_64_stage_1_0_t507;
reg [6-1:0] FSM_fft_64_stage_1_0_t508;
reg [64-1:0] FSM_fft_64_stage_1_0_t509;
reg [32-1:0] FSM_fft_64_stage_1_0_t510;
reg [6-1:0] FSM_fft_64_stage_1_0_t511;
reg [32-1:0] FSM_fft_64_stage_1_0_t512;
reg [64-1:0] FSM_fft_64_stage_1_0_t513;
reg [32-1:0] FSM_fft_64_stage_1_0_t514;
reg [33-1:0] FSM_fft_64_stage_1_0_t515;
reg [32-1:0] FSM_fft_64_stage_1_0_t516;
reg [6-1:0] FSM_fft_64_stage_1_0_t517;
reg [32-1:0] FSM_fft_64_stage_1_0_t518;
reg [33-1:0] FSM_fft_64_stage_1_0_t519;
reg [32-1:0] FSM_fft_64_stage_1_0_t520;
reg [2048-1:0] FSM_fft_64_stage_1_0_t521;
reg [64-1:0] FSM_fft_64_stage_1_0_t522;
reg [32-1:0] FSM_fft_64_stage_1_0_t523;
reg [33-1:0] FSM_fft_64_stage_1_0_t524;
reg [32-1:0] FSM_fft_64_stage_1_0_t525;
reg [6-1:0] FSM_fft_64_stage_1_0_t526;
reg [2048-1:0] FSM_fft_64_stage_1_0_t527;
reg [64-1:0] FSM_fft_64_stage_1_0_t528;
reg [32-1:0] FSM_fft_64_stage_1_0_t529;
reg [6-1:0] FSM_fft_64_stage_1_0_t530;
reg [64-1:0] FSM_fft_64_stage_1_0_t531;
reg [32-1:0] FSM_fft_64_stage_1_0_t532;
reg [6-1:0] FSM_fft_64_stage_1_0_t533;
reg [32-1:0] FSM_fft_64_stage_1_0_t534;
reg [64-1:0] FSM_fft_64_stage_1_0_t535;
reg [32-1:0] FSM_fft_64_stage_1_0_t536;
reg [33-1:0] FSM_fft_64_stage_1_0_t537;
reg [32-1:0] FSM_fft_64_stage_1_0_t538;
reg [6-1:0] FSM_fft_64_stage_1_0_t539;
reg [32-1:0] FSM_fft_64_stage_1_0_t540;
reg [33-1:0] FSM_fft_64_stage_1_0_t541;
reg [32-1:0] FSM_fft_64_stage_1_0_t542;
reg [2048-1:0] FSM_fft_64_stage_1_0_t543;
reg [64-1:0] FSM_fft_64_stage_1_0_t544;
reg [32-1:0] FSM_fft_64_stage_1_0_t545;
reg [33-1:0] FSM_fft_64_stage_1_0_t546;
reg [32-1:0] FSM_fft_64_stage_1_0_t547;
reg [6-1:0] FSM_fft_64_stage_1_0_t548;
reg [2048-1:0] FSM_fft_64_stage_1_0_t549;
reg [64-1:0] FSM_fft_64_stage_1_0_t550;
reg [32-1:0] FSM_fft_64_stage_1_0_t551;
reg [6-1:0] FSM_fft_64_stage_1_0_t552;
reg [64-1:0] FSM_fft_64_stage_1_0_t553;
reg [32-1:0] FSM_fft_64_stage_1_0_t554;
reg [6-1:0] FSM_fft_64_stage_1_0_t555;
reg [32-1:0] FSM_fft_64_stage_1_0_t556;
reg [64-1:0] FSM_fft_64_stage_1_0_t557;
reg [32-1:0] FSM_fft_64_stage_1_0_t558;
reg [33-1:0] FSM_fft_64_stage_1_0_t559;
reg [32-1:0] FSM_fft_64_stage_1_0_t560;
reg [6-1:0] FSM_fft_64_stage_1_0_t561;
reg [32-1:0] FSM_fft_64_stage_1_0_t562;
reg [33-1:0] FSM_fft_64_stage_1_0_t563;
reg [32-1:0] FSM_fft_64_stage_1_0_t564;
reg [2048-1:0] FSM_fft_64_stage_1_0_t565;
reg [64-1:0] FSM_fft_64_stage_1_0_t566;
reg [32-1:0] FSM_fft_64_stage_1_0_t567;
reg [33-1:0] FSM_fft_64_stage_1_0_t568;
reg [32-1:0] FSM_fft_64_stage_1_0_t569;
reg [6-1:0] FSM_fft_64_stage_1_0_t570;
reg [2048-1:0] FSM_fft_64_stage_1_0_t571;
reg [64-1:0] FSM_fft_64_stage_1_0_t572;
reg [32-1:0] FSM_fft_64_stage_1_0_t573;
reg [6-1:0] FSM_fft_64_stage_1_0_t574;
reg [64-1:0] FSM_fft_64_stage_1_0_t575;
reg [32-1:0] FSM_fft_64_stage_1_0_t576;
reg [6-1:0] FSM_fft_64_stage_1_0_t577;
reg [32-1:0] FSM_fft_64_stage_1_0_t578;
reg [64-1:0] FSM_fft_64_stage_1_0_t579;
reg [32-1:0] FSM_fft_64_stage_1_0_t580;
reg [33-1:0] FSM_fft_64_stage_1_0_t581;
reg [32-1:0] FSM_fft_64_stage_1_0_t582;
reg [6-1:0] FSM_fft_64_stage_1_0_t583;
reg [32-1:0] FSM_fft_64_stage_1_0_t584;
reg [33-1:0] FSM_fft_64_stage_1_0_t585;
reg [32-1:0] FSM_fft_64_stage_1_0_t586;
reg [2048-1:0] FSM_fft_64_stage_1_0_t587;
reg [64-1:0] FSM_fft_64_stage_1_0_t588;
reg [32-1:0] FSM_fft_64_stage_1_0_t589;
reg [33-1:0] FSM_fft_64_stage_1_0_t590;
reg [32-1:0] FSM_fft_64_stage_1_0_t591;
reg [6-1:0] FSM_fft_64_stage_1_0_t592;
reg [2048-1:0] FSM_fft_64_stage_1_0_t593;
reg [64-1:0] FSM_fft_64_stage_1_0_t594;
reg [32-1:0] FSM_fft_64_stage_1_0_t595;
reg [6-1:0] FSM_fft_64_stage_1_0_t596;
reg [64-1:0] FSM_fft_64_stage_1_0_t597;
reg [32-1:0] FSM_fft_64_stage_1_0_t598;
reg [6-1:0] FSM_fft_64_stage_1_0_t599;
reg [32-1:0] FSM_fft_64_stage_1_0_t600;
reg [64-1:0] FSM_fft_64_stage_1_0_t601;
reg [32-1:0] FSM_fft_64_stage_1_0_t602;
reg [33-1:0] FSM_fft_64_stage_1_0_t603;
reg [32-1:0] FSM_fft_64_stage_1_0_t604;
reg [6-1:0] FSM_fft_64_stage_1_0_t605;
reg [32-1:0] FSM_fft_64_stage_1_0_t606;
reg [33-1:0] FSM_fft_64_stage_1_0_t607;
reg [32-1:0] FSM_fft_64_stage_1_0_t608;
reg [2048-1:0] FSM_fft_64_stage_1_0_t609;
reg [64-1:0] FSM_fft_64_stage_1_0_t610;
reg [32-1:0] FSM_fft_64_stage_1_0_t611;
reg [33-1:0] FSM_fft_64_stage_1_0_t612;
reg [32-1:0] FSM_fft_64_stage_1_0_t613;
reg [6-1:0] FSM_fft_64_stage_1_0_t614;
reg [2048-1:0] FSM_fft_64_stage_1_0_t615;
reg [64-1:0] FSM_fft_64_stage_1_0_t616;
reg [32-1:0] FSM_fft_64_stage_1_0_t617;
reg [6-1:0] FSM_fft_64_stage_1_0_t618;
reg [64-1:0] FSM_fft_64_stage_1_0_t619;
reg [32-1:0] FSM_fft_64_stage_1_0_t620;
reg [6-1:0] FSM_fft_64_stage_1_0_t621;
reg [32-1:0] FSM_fft_64_stage_1_0_t622;
reg [64-1:0] FSM_fft_64_stage_1_0_t623;
reg [32-1:0] FSM_fft_64_stage_1_0_t624;
reg [33-1:0] FSM_fft_64_stage_1_0_t625;
reg [32-1:0] FSM_fft_64_stage_1_0_t626;
reg [6-1:0] FSM_fft_64_stage_1_0_t627;
reg [32-1:0] FSM_fft_64_stage_1_0_t628;
reg [33-1:0] FSM_fft_64_stage_1_0_t629;
reg [32-1:0] FSM_fft_64_stage_1_0_t630;
reg [2048-1:0] FSM_fft_64_stage_1_0_t631;
reg [64-1:0] FSM_fft_64_stage_1_0_t632;
reg [32-1:0] FSM_fft_64_stage_1_0_t633;
reg [33-1:0] FSM_fft_64_stage_1_0_t634;
reg [32-1:0] FSM_fft_64_stage_1_0_t635;
reg [6-1:0] FSM_fft_64_stage_1_0_t636;
reg [2048-1:0] FSM_fft_64_stage_1_0_t637;
reg [64-1:0] FSM_fft_64_stage_1_0_t638;
reg [32-1:0] FSM_fft_64_stage_1_0_t639;
reg [6-1:0] FSM_fft_64_stage_1_0_t640;
reg [64-1:0] FSM_fft_64_stage_1_0_t641;
reg [32-1:0] FSM_fft_64_stage_1_0_t642;
reg [6-1:0] FSM_fft_64_stage_1_0_t643;
reg [32-1:0] FSM_fft_64_stage_1_0_t644;
reg [64-1:0] FSM_fft_64_stage_1_0_t645;
reg [32-1:0] FSM_fft_64_stage_1_0_t646;
reg [33-1:0] FSM_fft_64_stage_1_0_t647;
reg [32-1:0] FSM_fft_64_stage_1_0_t648;
reg [6-1:0] FSM_fft_64_stage_1_0_t649;
reg [32-1:0] FSM_fft_64_stage_1_0_t650;
reg [33-1:0] FSM_fft_64_stage_1_0_t651;
reg [32-1:0] FSM_fft_64_stage_1_0_t652;
reg [2048-1:0] FSM_fft_64_stage_1_0_t653;
reg [64-1:0] FSM_fft_64_stage_1_0_t654;
reg [32-1:0] FSM_fft_64_stage_1_0_t655;
reg [33-1:0] FSM_fft_64_stage_1_0_t656;
reg [32-1:0] FSM_fft_64_stage_1_0_t657;
reg [6-1:0] FSM_fft_64_stage_1_0_t658;
reg [2048-1:0] FSM_fft_64_stage_1_0_t659;
reg [64-1:0] FSM_fft_64_stage_1_0_t660;
reg [32-1:0] FSM_fft_64_stage_1_0_t661;
reg [6-1:0] FSM_fft_64_stage_1_0_t662;
reg [64-1:0] FSM_fft_64_stage_1_0_t663;
reg [32-1:0] FSM_fft_64_stage_1_0_t664;
reg [6-1:0] FSM_fft_64_stage_1_0_t665;
reg [32-1:0] FSM_fft_64_stage_1_0_t666;
reg [64-1:0] FSM_fft_64_stage_1_0_t667;
reg [32-1:0] FSM_fft_64_stage_1_0_t668;
reg [33-1:0] FSM_fft_64_stage_1_0_t669;
reg [32-1:0] FSM_fft_64_stage_1_0_t670;
reg [6-1:0] FSM_fft_64_stage_1_0_t671;
reg [32-1:0] FSM_fft_64_stage_1_0_t672;
reg [33-1:0] FSM_fft_64_stage_1_0_t673;
reg [32-1:0] FSM_fft_64_stage_1_0_t674;
reg [2048-1:0] FSM_fft_64_stage_1_0_t675;
reg [64-1:0] FSM_fft_64_stage_1_0_t676;
reg [32-1:0] FSM_fft_64_stage_1_0_t677;
reg [33-1:0] FSM_fft_64_stage_1_0_t678;
reg [32-1:0] FSM_fft_64_stage_1_0_t679;
reg [6-1:0] FSM_fft_64_stage_1_0_t680;
reg [2048-1:0] FSM_fft_64_stage_1_0_t681;
reg [64-1:0] FSM_fft_64_stage_1_0_t682;
reg [32-1:0] FSM_fft_64_stage_1_0_t683;
reg [6-1:0] FSM_fft_64_stage_1_0_t684;
reg [64-1:0] FSM_fft_64_stage_1_0_t685;
reg [32-1:0] FSM_fft_64_stage_1_0_t686;
reg [6-1:0] FSM_fft_64_stage_1_0_t687;
reg [32-1:0] FSM_fft_64_stage_1_0_t688;
reg [64-1:0] FSM_fft_64_stage_1_0_t689;
reg [32-1:0] FSM_fft_64_stage_1_0_t690;
reg [33-1:0] FSM_fft_64_stage_1_0_t691;
reg [32-1:0] FSM_fft_64_stage_1_0_t692;
reg [6-1:0] FSM_fft_64_stage_1_0_t693;
reg [32-1:0] FSM_fft_64_stage_1_0_t694;
reg [33-1:0] FSM_fft_64_stage_1_0_t695;
reg [32-1:0] FSM_fft_64_stage_1_0_t696;
reg [2048-1:0] FSM_fft_64_stage_1_0_t697;
reg [64-1:0] FSM_fft_64_stage_1_0_t698;
reg [32-1:0] FSM_fft_64_stage_1_0_t699;
reg [33-1:0] FSM_fft_64_stage_1_0_t700;
reg [32-1:0] FSM_fft_64_stage_1_0_t701;
reg [6-1:0] FSM_fft_64_stage_1_0_t702;
reg [2048-1:0] FSM_fft_64_stage_1_0_t703;
reg [64-1:0] FSM_fft_64_stage_1_0_t704;
reg [32-1:0] FSM_fft_64_stage_1_0_t705;
reg [6-1:0] FSM_fft_64_stage_1_0_t706;
reg [64-1:0] FSM_fft_64_stage_1_0_t707;
reg [32-1:0] FSM_fft_64_stage_1_0_t708;
reg [6-1:0] FSM_fft_64_stage_1_0_t709;
reg [32-1:0] FSM_fft_64_stage_1_0_t710;
reg [64-1:0] FSM_fft_64_stage_1_0_t711;
reg [32-1:0] FSM_fft_64_stage_1_0_t712;
reg [33-1:0] FSM_fft_64_stage_1_0_t713;
reg [32-1:0] FSM_fft_64_stage_1_0_t714;
reg [6-1:0] FSM_fft_64_stage_1_0_t715;
reg [32-1:0] FSM_fft_64_stage_1_0_t716;
reg [33-1:0] FSM_fft_64_stage_1_0_t717;
reg [32-1:0] FSM_fft_64_stage_1_0_t718;
reg [2048-1:0] FSM_fft_64_stage_1_0_t719;
reg [64-1:0] FSM_fft_64_stage_1_0_t720;
reg [32-1:0] FSM_fft_64_stage_1_0_t721;
reg [33-1:0] FSM_fft_64_stage_1_0_t722;
reg [32-1:0] FSM_fft_64_stage_1_0_t723;
reg [6-1:0] FSM_fft_64_stage_1_0_t724;
reg [2048-1:0] FSM_fft_64_stage_1_0_t725;
reg [64-1:0] FSM_fft_64_stage_1_0_t726;
reg [32-1:0] FSM_fft_64_stage_1_0_t727;
reg [6-1:0] FSM_fft_64_stage_1_0_t728;
reg [64-1:0] FSM_fft_64_stage_1_0_t729;
reg [32-1:0] FSM_fft_64_stage_1_0_t730;
reg [6-1:0] FSM_fft_64_stage_1_0_t731;
reg [32-1:0] FSM_fft_64_stage_1_0_t732;
reg [64-1:0] FSM_fft_64_stage_1_0_t733;
reg [32-1:0] FSM_fft_64_stage_1_0_t734;
reg [33-1:0] FSM_fft_64_stage_1_0_t735;
reg [32-1:0] FSM_fft_64_stage_1_0_t736;
reg [6-1:0] FSM_fft_64_stage_1_0_t737;
reg [32-1:0] FSM_fft_64_stage_1_0_t738;
reg [33-1:0] FSM_fft_64_stage_1_0_t739;
reg [32-1:0] FSM_fft_64_stage_1_0_t740;
reg [2048-1:0] FSM_fft_64_stage_1_0_t741;
reg [64-1:0] FSM_fft_64_stage_1_0_t742;
reg [32-1:0] FSM_fft_64_stage_1_0_t743;
reg [33-1:0] FSM_fft_64_stage_1_0_t744;
reg [32-1:0] FSM_fft_64_stage_1_0_t745;
reg [6-1:0] FSM_fft_64_stage_1_0_t746;
reg [2048-1:0] FSM_fft_64_stage_1_0_t747;
reg [64-1:0] FSM_fft_64_stage_1_0_t748;
reg [32-1:0] FSM_fft_64_stage_1_0_t749;
reg [6-1:0] FSM_fft_64_stage_1_0_t750;
reg [64-1:0] FSM_fft_64_stage_1_0_t751;
reg [32-1:0] FSM_fft_64_stage_1_0_t752;
reg [6-1:0] FSM_fft_64_stage_1_0_t753;
reg [32-1:0] FSM_fft_64_stage_1_0_t754;
reg [64-1:0] FSM_fft_64_stage_1_0_t755;
reg [32-1:0] FSM_fft_64_stage_1_0_t756;
reg [33-1:0] FSM_fft_64_stage_1_0_t757;
reg [32-1:0] FSM_fft_64_stage_1_0_t758;
reg [6-1:0] FSM_fft_64_stage_1_0_t759;
reg [32-1:0] FSM_fft_64_stage_1_0_t760;
reg [33-1:0] FSM_fft_64_stage_1_0_t761;
reg [32-1:0] FSM_fft_64_stage_1_0_t762;
reg [2048-1:0] FSM_fft_64_stage_1_0_t763;
reg [64-1:0] FSM_fft_64_stage_1_0_t764;
reg [32-1:0] FSM_fft_64_stage_1_0_t765;
reg [33-1:0] FSM_fft_64_stage_1_0_t766;
reg [32-1:0] FSM_fft_64_stage_1_0_t767;
reg [6-1:0] FSM_fft_64_stage_1_0_t768;
reg [2048-1:0] FSM_fft_64_stage_1_0_t769;
reg [64-1:0] FSM_fft_64_stage_1_0_t770;
reg [32-1:0] FSM_fft_64_stage_1_0_t771;
reg [6-1:0] FSM_fft_64_stage_1_0_t772;
reg [64-1:0] FSM_fft_64_stage_1_0_t773;
reg [32-1:0] FSM_fft_64_stage_1_0_t774;
reg [6-1:0] FSM_fft_64_stage_1_0_t775;
reg [32-1:0] FSM_fft_64_stage_1_0_t776;
reg [64-1:0] FSM_fft_64_stage_1_0_t777;
reg [32-1:0] FSM_fft_64_stage_1_0_t778;
reg [33-1:0] FSM_fft_64_stage_1_0_t779;
reg [32-1:0] FSM_fft_64_stage_1_0_t780;
reg [6-1:0] FSM_fft_64_stage_1_0_t781;
reg [32-1:0] FSM_fft_64_stage_1_0_t782;
reg [33-1:0] FSM_fft_64_stage_1_0_t783;
reg [32-1:0] FSM_fft_64_stage_1_0_t784;
reg [2048-1:0] FSM_fft_64_stage_1_0_t785;
reg [64-1:0] FSM_fft_64_stage_1_0_t786;
reg [32-1:0] FSM_fft_64_stage_1_0_t787;
reg [33-1:0] FSM_fft_64_stage_1_0_t788;
reg [32-1:0] FSM_fft_64_stage_1_0_t789;
reg [6-1:0] FSM_fft_64_stage_1_0_t790;
reg [2048-1:0] FSM_fft_64_stage_1_0_t791;
reg [64-1:0] FSM_fft_64_stage_1_0_t792;
reg [32-1:0] FSM_fft_64_stage_1_0_t793;
reg [6-1:0] FSM_fft_64_stage_1_0_t794;
reg [64-1:0] FSM_fft_64_stage_1_0_t795;
reg [32-1:0] FSM_fft_64_stage_1_0_t796;
reg [6-1:0] FSM_fft_64_stage_1_0_t797;
reg [32-1:0] FSM_fft_64_stage_1_0_t798;
reg [64-1:0] FSM_fft_64_stage_1_0_t799;
reg [32-1:0] FSM_fft_64_stage_1_0_t800;
reg [33-1:0] FSM_fft_64_stage_1_0_t801;
reg [32-1:0] FSM_fft_64_stage_1_0_t802;
reg [6-1:0] FSM_fft_64_stage_1_0_t803;
reg [32-1:0] FSM_fft_64_stage_1_0_t804;
reg [33-1:0] FSM_fft_64_stage_1_0_t805;
reg [32-1:0] FSM_fft_64_stage_1_0_t806;
reg [2048-1:0] FSM_fft_64_stage_1_0_t807;
reg [64-1:0] FSM_fft_64_stage_1_0_t808;
reg [32-1:0] FSM_fft_64_stage_1_0_t809;
reg [33-1:0] FSM_fft_64_stage_1_0_t810;
reg [32-1:0] FSM_fft_64_stage_1_0_t811;
reg [6-1:0] FSM_fft_64_stage_1_0_t812;
reg [2048-1:0] FSM_fft_64_stage_1_0_t813;
reg [64-1:0] FSM_fft_64_stage_1_0_t814;
reg [32-1:0] FSM_fft_64_stage_1_0_t815;
reg [6-1:0] FSM_fft_64_stage_1_0_t816;
reg [64-1:0] FSM_fft_64_stage_1_0_t817;
reg [32-1:0] FSM_fft_64_stage_1_0_t818;
reg [6-1:0] FSM_fft_64_stage_1_0_t819;
reg [32-1:0] FSM_fft_64_stage_1_0_t820;
reg [64-1:0] FSM_fft_64_stage_1_0_t821;
reg [32-1:0] FSM_fft_64_stage_1_0_t822;
reg [33-1:0] FSM_fft_64_stage_1_0_t823;
reg [32-1:0] FSM_fft_64_stage_1_0_t824;
reg [6-1:0] FSM_fft_64_stage_1_0_t825;
reg [32-1:0] FSM_fft_64_stage_1_0_t826;
reg [33-1:0] FSM_fft_64_stage_1_0_t827;
reg [32-1:0] FSM_fft_64_stage_1_0_t828;
reg [2048-1:0] FSM_fft_64_stage_1_0_t829;
reg [64-1:0] FSM_fft_64_stage_1_0_t830;
reg [32-1:0] FSM_fft_64_stage_1_0_t831;
reg [33-1:0] FSM_fft_64_stage_1_0_t832;
reg [32-1:0] FSM_fft_64_stage_1_0_t833;
reg [6-1:0] FSM_fft_64_stage_1_0_t834;
reg [2048-1:0] FSM_fft_64_stage_1_0_t835;
reg [64-1:0] FSM_fft_64_stage_1_0_t836;
reg [32-1:0] FSM_fft_64_stage_1_0_t837;
reg [6-1:0] FSM_fft_64_stage_1_0_t838;
reg [64-1:0] FSM_fft_64_stage_1_0_t839;
reg [32-1:0] FSM_fft_64_stage_1_0_t840;
reg [6-1:0] FSM_fft_64_stage_1_0_t841;
reg [32-1:0] FSM_fft_64_stage_1_0_t842;
reg [64-1:0] FSM_fft_64_stage_1_0_t843;
reg [32-1:0] FSM_fft_64_stage_1_0_t844;
reg [33-1:0] FSM_fft_64_stage_1_0_t845;
reg [32-1:0] FSM_fft_64_stage_1_0_t846;
reg [6-1:0] FSM_fft_64_stage_1_0_t847;
reg [32-1:0] FSM_fft_64_stage_1_0_t848;
reg [33-1:0] FSM_fft_64_stage_1_0_t849;
reg [32-1:0] FSM_fft_64_stage_1_0_t850;
reg [2048-1:0] FSM_fft_64_stage_1_0_t851;
reg [64-1:0] FSM_fft_64_stage_1_0_t852;
reg [32-1:0] FSM_fft_64_stage_1_0_t853;
reg [33-1:0] FSM_fft_64_stage_1_0_t854;
reg [32-1:0] FSM_fft_64_stage_1_0_t855;
reg [6-1:0] FSM_fft_64_stage_1_0_t856;
reg [2048-1:0] FSM_fft_64_stage_1_0_t857;
reg [64-1:0] FSM_fft_64_stage_1_0_t858;
reg [32-1:0] FSM_fft_64_stage_1_0_t859;
reg [6-1:0] FSM_fft_64_stage_1_0_t860;
reg [64-1:0] FSM_fft_64_stage_1_0_t861;
reg [32-1:0] FSM_fft_64_stage_1_0_t862;
reg [6-1:0] FSM_fft_64_stage_1_0_t863;
reg [32-1:0] FSM_fft_64_stage_1_0_t864;
reg [64-1:0] FSM_fft_64_stage_1_0_t865;
reg [32-1:0] FSM_fft_64_stage_1_0_t866;
reg [33-1:0] FSM_fft_64_stage_1_0_t867;
reg [32-1:0] FSM_fft_64_stage_1_0_t868;
reg [6-1:0] FSM_fft_64_stage_1_0_t869;
reg [32-1:0] FSM_fft_64_stage_1_0_t870;
reg [33-1:0] FSM_fft_64_stage_1_0_t871;
reg [32-1:0] FSM_fft_64_stage_1_0_t872;
reg [2048-1:0] FSM_fft_64_stage_1_0_t873;
reg [64-1:0] FSM_fft_64_stage_1_0_t874;
reg [32-1:0] FSM_fft_64_stage_1_0_t875;
reg [33-1:0] FSM_fft_64_stage_1_0_t876;
reg [32-1:0] FSM_fft_64_stage_1_0_t877;
reg [6-1:0] FSM_fft_64_stage_1_0_t878;
reg [2048-1:0] FSM_fft_64_stage_1_0_t879;
reg [64-1:0] FSM_fft_64_stage_1_0_t880;
reg [32-1:0] FSM_fft_64_stage_1_0_t881;
reg [6-1:0] FSM_fft_64_stage_1_0_t882;
reg [64-1:0] FSM_fft_64_stage_1_0_t883;
reg [32-1:0] FSM_fft_64_stage_1_0_t884;
reg [6-1:0] FSM_fft_64_stage_1_0_t885;
reg [32-1:0] FSM_fft_64_stage_1_0_t886;
reg [64-1:0] FSM_fft_64_stage_1_0_t887;
reg [32-1:0] FSM_fft_64_stage_1_0_t888;
reg [33-1:0] FSM_fft_64_stage_1_0_t889;
reg [32-1:0] FSM_fft_64_stage_1_0_t890;
reg [6-1:0] FSM_fft_64_stage_1_0_t891;
reg [32-1:0] FSM_fft_64_stage_1_0_t892;
reg [33-1:0] FSM_fft_64_stage_1_0_t893;
reg [32-1:0] FSM_fft_64_stage_1_0_t894;
reg [2048-1:0] FSM_fft_64_stage_1_0_t895;
reg [64-1:0] FSM_fft_64_stage_1_0_t896;
reg [32-1:0] FSM_fft_64_stage_1_0_t897;
reg [33-1:0] FSM_fft_64_stage_1_0_t898;
reg [32-1:0] FSM_fft_64_stage_1_0_t899;
reg [6-1:0] FSM_fft_64_stage_1_0_t900;
reg [2048-1:0] FSM_fft_64_stage_1_0_t901;
reg [64-1:0] FSM_fft_64_stage_1_0_t902;
reg [32-1:0] FSM_fft_64_stage_1_0_t903;
reg [6-1:0] FSM_fft_64_stage_1_0_t904;
reg [64-1:0] FSM_fft_64_stage_1_0_t905;
reg [32-1:0] FSM_fft_64_stage_1_0_t906;
reg [6-1:0] FSM_fft_64_stage_1_0_t907;
reg [32-1:0] FSM_fft_64_stage_1_0_t908;
reg [64-1:0] FSM_fft_64_stage_1_0_t909;
reg [32-1:0] FSM_fft_64_stage_1_0_t910;
reg [33-1:0] FSM_fft_64_stage_1_0_t911;
reg [32-1:0] FSM_fft_64_stage_1_0_t912;
reg [6-1:0] FSM_fft_64_stage_1_0_t913;
reg [32-1:0] FSM_fft_64_stage_1_0_t914;
reg [33-1:0] FSM_fft_64_stage_1_0_t915;
reg [32-1:0] FSM_fft_64_stage_1_0_t916;
reg [2048-1:0] FSM_fft_64_stage_1_0_t917;
reg [64-1:0] FSM_fft_64_stage_1_0_t918;
reg [32-1:0] FSM_fft_64_stage_1_0_t919;
reg [33-1:0] FSM_fft_64_stage_1_0_t920;
reg [32-1:0] FSM_fft_64_stage_1_0_t921;
reg [6-1:0] FSM_fft_64_stage_1_0_t922;
reg [2048-1:0] FSM_fft_64_stage_1_0_t923;
reg [64-1:0] FSM_fft_64_stage_1_0_t924;
reg [32-1:0] FSM_fft_64_stage_1_0_t925;
reg [6-1:0] FSM_fft_64_stage_1_0_t926;
reg [64-1:0] FSM_fft_64_stage_1_0_t927;
reg [32-1:0] FSM_fft_64_stage_1_0_t928;
reg [6-1:0] FSM_fft_64_stage_1_0_t929;
reg [32-1:0] FSM_fft_64_stage_1_0_t930;
reg [64-1:0] FSM_fft_64_stage_1_0_t931;
reg [32-1:0] FSM_fft_64_stage_1_0_t932;
reg [33-1:0] FSM_fft_64_stage_1_0_t933;
reg [32-1:0] FSM_fft_64_stage_1_0_t934;
reg [6-1:0] FSM_fft_64_stage_1_0_t935;
reg [32-1:0] FSM_fft_64_stage_1_0_t936;
reg [33-1:0] FSM_fft_64_stage_1_0_t937;
reg [32-1:0] FSM_fft_64_stage_1_0_t938;
reg [2048-1:0] FSM_fft_64_stage_1_0_t939;
reg [64-1:0] FSM_fft_64_stage_1_0_t940;
reg [32-1:0] FSM_fft_64_stage_1_0_t941;
reg [33-1:0] FSM_fft_64_stage_1_0_t942;
reg [32-1:0] FSM_fft_64_stage_1_0_t943;
reg [6-1:0] FSM_fft_64_stage_1_0_t944;
reg [2048-1:0] FSM_fft_64_stage_1_0_t945;
reg [64-1:0] FSM_fft_64_stage_1_0_t946;
reg [32-1:0] FSM_fft_64_stage_1_0_t947;
reg [6-1:0] FSM_fft_64_stage_1_0_t948;
reg [64-1:0] FSM_fft_64_stage_1_0_t949;
reg [32-1:0] FSM_fft_64_stage_1_0_t950;
reg [6-1:0] FSM_fft_64_stage_1_0_t951;
reg [32-1:0] FSM_fft_64_stage_1_0_t952;
reg [64-1:0] FSM_fft_64_stage_1_0_t953;
reg [32-1:0] FSM_fft_64_stage_1_0_t954;
reg [33-1:0] FSM_fft_64_stage_1_0_t955;
reg [32-1:0] FSM_fft_64_stage_1_0_t956;
reg [6-1:0] FSM_fft_64_stage_1_0_t957;
reg [32-1:0] FSM_fft_64_stage_1_0_t958;
reg [33-1:0] FSM_fft_64_stage_1_0_t959;
reg [32-1:0] FSM_fft_64_stage_1_0_t960;
reg [2048-1:0] FSM_fft_64_stage_1_0_t961;
reg [64-1:0] FSM_fft_64_stage_1_0_t962;
reg [32-1:0] FSM_fft_64_stage_1_0_t963;
reg [33-1:0] FSM_fft_64_stage_1_0_t964;
reg [32-1:0] FSM_fft_64_stage_1_0_t965;
reg [6-1:0] FSM_fft_64_stage_1_0_t966;
reg [2048-1:0] FSM_fft_64_stage_1_0_t967;
reg [64-1:0] FSM_fft_64_stage_1_0_t968;
reg [32-1:0] FSM_fft_64_stage_1_0_t969;
reg [6-1:0] FSM_fft_64_stage_1_0_t970;
reg [64-1:0] FSM_fft_64_stage_1_0_t971;
reg [32-1:0] FSM_fft_64_stage_1_0_t972;
reg [6-1:0] FSM_fft_64_stage_1_0_t973;
reg [32-1:0] FSM_fft_64_stage_1_0_t974;
reg [64-1:0] FSM_fft_64_stage_1_0_t975;
reg [32-1:0] FSM_fft_64_stage_1_0_t976;
reg [33-1:0] FSM_fft_64_stage_1_0_t977;
reg [32-1:0] FSM_fft_64_stage_1_0_t978;
reg [6-1:0] FSM_fft_64_stage_1_0_t979;
reg [32-1:0] FSM_fft_64_stage_1_0_t980;
reg [33-1:0] FSM_fft_64_stage_1_0_t981;
reg [32-1:0] FSM_fft_64_stage_1_0_t982;
reg [2048-1:0] FSM_fft_64_stage_1_0_t983;
reg [64-1:0] FSM_fft_64_stage_1_0_t984;
reg [32-1:0] FSM_fft_64_stage_1_0_t985;
reg [33-1:0] FSM_fft_64_stage_1_0_t986;
reg [32-1:0] FSM_fft_64_stage_1_0_t987;
reg [6-1:0] FSM_fft_64_stage_1_0_t988;
reg [2048-1:0] FSM_fft_64_stage_1_0_t989;
reg [64-1:0] FSM_fft_64_stage_1_0_t990;
reg [32-1:0] FSM_fft_64_stage_1_0_t991;
reg [6-1:0] FSM_fft_64_stage_1_0_t992;
reg [64-1:0] FSM_fft_64_stage_1_0_t993;
reg [32-1:0] FSM_fft_64_stage_1_0_t994;
reg [6-1:0] FSM_fft_64_stage_1_0_t995;
reg [32-1:0] FSM_fft_64_stage_1_0_t996;
reg [64-1:0] FSM_fft_64_stage_1_0_t997;
reg [32-1:0] FSM_fft_64_stage_1_0_t998;
reg [33-1:0] FSM_fft_64_stage_1_0_t999;
reg [32-1:0] FSM_fft_64_stage_1_0_t1000;
reg [6-1:0] FSM_fft_64_stage_1_0_t1001;
reg [32-1:0] FSM_fft_64_stage_1_0_t1002;
reg [33-1:0] FSM_fft_64_stage_1_0_t1003;
reg [32-1:0] FSM_fft_64_stage_1_0_t1004;
reg [2048-1:0] FSM_fft_64_stage_1_0_t1005;
reg [64-1:0] FSM_fft_64_stage_1_0_t1006;
reg [32-1:0] FSM_fft_64_stage_1_0_t1007;
reg [33-1:0] FSM_fft_64_stage_1_0_t1008;
reg [32-1:0] FSM_fft_64_stage_1_0_t1009;
reg [6-1:0] FSM_fft_64_stage_1_0_t1010;
reg [2048-1:0] FSM_fft_64_stage_1_0_t1011;
reg [64-1:0] FSM_fft_64_stage_1_0_t1012;
reg [32-1:0] FSM_fft_64_stage_1_0_t1013;
reg [6-1:0] FSM_fft_64_stage_1_0_t1014;
reg [64-1:0] FSM_fft_64_stage_1_0_t1015;
reg [32-1:0] FSM_fft_64_stage_1_0_t1016;
reg [6-1:0] FSM_fft_64_stage_1_0_t1017;
reg [32-1:0] FSM_fft_64_stage_1_0_t1018;
reg [64-1:0] FSM_fft_64_stage_1_0_t1019;
reg [32-1:0] FSM_fft_64_stage_1_0_t1020;
reg [33-1:0] FSM_fft_64_stage_1_0_t1021;
reg [32-1:0] FSM_fft_64_stage_1_0_t1022;
reg [6-1:0] FSM_fft_64_stage_1_0_t1023;
reg [32-1:0] FSM_fft_64_stage_1_0_t1024;
reg [33-1:0] FSM_fft_64_stage_1_0_t1025;
reg [32-1:0] FSM_fft_64_stage_1_0_t1026;
reg [2048-1:0] FSM_fft_64_stage_1_0_t1027;
reg [64-1:0] FSM_fft_64_stage_1_0_t1028;
reg [32-1:0] FSM_fft_64_stage_1_0_t1029;
reg [33-1:0] FSM_fft_64_stage_1_0_t1030;
reg [32-1:0] FSM_fft_64_stage_1_0_t1031;
reg [6-1:0] FSM_fft_64_stage_1_0_t1032;
reg [2048-1:0] FSM_fft_64_stage_1_0_t1033;
reg [64-1:0] FSM_fft_64_stage_1_0_t1034;
reg [32-1:0] FSM_fft_64_stage_1_0_t1035;
reg [6-1:0] FSM_fft_64_stage_1_0_t1036;
reg [64-1:0] FSM_fft_64_stage_1_0_t1037;
reg [32-1:0] FSM_fft_64_stage_1_0_t1038;
reg [6-1:0] FSM_fft_64_stage_1_0_t1039;
reg [32-1:0] FSM_fft_64_stage_1_0_t1040;
reg [64-1:0] FSM_fft_64_stage_1_0_t1041;
reg [32-1:0] FSM_fft_64_stage_1_0_t1042;
reg [33-1:0] FSM_fft_64_stage_1_0_t1043;
reg [32-1:0] FSM_fft_64_stage_1_0_t1044;
reg [6-1:0] FSM_fft_64_stage_1_0_t1045;
reg [32-1:0] FSM_fft_64_stage_1_0_t1046;
reg [33-1:0] FSM_fft_64_stage_1_0_t1047;
reg [32-1:0] FSM_fft_64_stage_1_0_t1048;
reg [2048-1:0] FSM_fft_64_stage_1_0_t1049;
reg [64-1:0] FSM_fft_64_stage_1_0_t1050;
reg [32-1:0] FSM_fft_64_stage_1_0_t1051;
reg [33-1:0] FSM_fft_64_stage_1_0_t1052;
reg [32-1:0] FSM_fft_64_stage_1_0_t1053;
reg [6-1:0] FSM_fft_64_stage_1_0_t1054;
reg [2048-1:0] FSM_fft_64_stage_1_0_t1055;
reg [64-1:0] FSM_fft_64_stage_1_0_t1056;
reg [32-1:0] FSM_fft_64_stage_1_0_t1057;
reg [6-1:0] FSM_fft_64_stage_1_0_t1058;
reg [64-1:0] FSM_fft_64_stage_1_0_t1059;
reg [32-1:0] FSM_fft_64_stage_1_0_t1060;
reg [6-1:0] FSM_fft_64_stage_1_0_t1061;
reg [32-1:0] FSM_fft_64_stage_1_0_t1062;
reg [64-1:0] FSM_fft_64_stage_1_0_t1063;
reg [32-1:0] FSM_fft_64_stage_1_0_t1064;
reg [33-1:0] FSM_fft_64_stage_1_0_t1065;
reg [32-1:0] FSM_fft_64_stage_1_0_t1066;
reg [6-1:0] FSM_fft_64_stage_1_0_t1067;
reg [32-1:0] FSM_fft_64_stage_1_0_t1068;
reg [33-1:0] FSM_fft_64_stage_1_0_t1069;
reg [32-1:0] FSM_fft_64_stage_1_0_t1070;
reg [2048-1:0] FSM_fft_64_stage_1_0_t1071;
reg [64-1:0] FSM_fft_64_stage_1_0_t1072;
reg [32-1:0] FSM_fft_64_stage_1_0_t1073;
reg [33-1:0] FSM_fft_64_stage_1_0_t1074;
reg [32-1:0] FSM_fft_64_stage_1_0_t1075;
reg [6-1:0] FSM_fft_64_stage_1_0_t1076;
reg [2048-1:0] FSM_fft_64_stage_1_0_t1077;
reg [64-1:0] FSM_fft_64_stage_1_0_t1078;
reg [32-1:0] FSM_fft_64_stage_1_0_t1079;
reg [6-1:0] FSM_fft_64_stage_1_0_t1080;
reg [64-1:0] FSM_fft_64_stage_1_0_t1081;
reg [32-1:0] FSM_fft_64_stage_1_0_t1082;
reg [6-1:0] FSM_fft_64_stage_1_0_t1083;
reg [32-1:0] FSM_fft_64_stage_1_0_t1084;
reg [64-1:0] FSM_fft_64_stage_1_0_t1085;
reg [32-1:0] FSM_fft_64_stage_1_0_t1086;
reg [33-1:0] FSM_fft_64_stage_1_0_t1087;
reg [32-1:0] FSM_fft_64_stage_1_0_t1088;
reg [6-1:0] FSM_fft_64_stage_1_0_t1089;
reg [32-1:0] FSM_fft_64_stage_1_0_t1090;
reg [33-1:0] FSM_fft_64_stage_1_0_t1091;
reg [32-1:0] FSM_fft_64_stage_1_0_t1092;
reg [2048-1:0] FSM_fft_64_stage_1_0_t1093;
reg [64-1:0] FSM_fft_64_stage_1_0_t1094;
reg [32-1:0] FSM_fft_64_stage_1_0_t1095;
reg [33-1:0] FSM_fft_64_stage_1_0_t1096;
reg [32-1:0] FSM_fft_64_stage_1_0_t1097;
reg [6-1:0] FSM_fft_64_stage_1_0_t1098;
reg [2048-1:0] FSM_fft_64_stage_1_0_t1099;
reg [64-1:0] FSM_fft_64_stage_1_0_t1100;
reg [32-1:0] FSM_fft_64_stage_1_0_t1101;
reg [6-1:0] FSM_fft_64_stage_1_0_t1102;
reg [64-1:0] FSM_fft_64_stage_1_0_t1103;
reg [32-1:0] FSM_fft_64_stage_1_0_t1104;
reg [6-1:0] FSM_fft_64_stage_1_0_t1105;
reg [32-1:0] FSM_fft_64_stage_1_0_t1106;
reg [64-1:0] FSM_fft_64_stage_1_0_t1107;
reg [32-1:0] FSM_fft_64_stage_1_0_t1108;
reg [33-1:0] FSM_fft_64_stage_1_0_t1109;
reg [32-1:0] FSM_fft_64_stage_1_0_t1110;
reg [6-1:0] FSM_fft_64_stage_1_0_t1111;
reg [32-1:0] FSM_fft_64_stage_1_0_t1112;
reg [33-1:0] FSM_fft_64_stage_1_0_t1113;
reg [32-1:0] FSM_fft_64_stage_1_0_t1114;
reg [2048-1:0] FSM_fft_64_stage_1_0_t1115;
reg [64-1:0] FSM_fft_64_stage_1_0_t1116;
reg [32-1:0] FSM_fft_64_stage_1_0_t1117;
reg [33-1:0] FSM_fft_64_stage_1_0_t1118;
reg [32-1:0] FSM_fft_64_stage_1_0_t1119;
reg [6-1:0] FSM_fft_64_stage_1_0_t1120;
reg [2048-1:0] FSM_fft_64_stage_1_0_t1121;
reg [64-1:0] FSM_fft_64_stage_1_0_t1122;
reg [32-1:0] FSM_fft_64_stage_1_0_t1123;
reg [6-1:0] FSM_fft_64_stage_1_0_t1124;
reg [64-1:0] FSM_fft_64_stage_1_0_t1125;
reg [32-1:0] FSM_fft_64_stage_1_0_t1126;
reg [6-1:0] FSM_fft_64_stage_1_0_t1127;
reg [32-1:0] FSM_fft_64_stage_1_0_t1128;
reg [64-1:0] FSM_fft_64_stage_1_0_t1129;
reg [32-1:0] FSM_fft_64_stage_1_0_t1130;
reg [33-1:0] FSM_fft_64_stage_1_0_t1131;
reg [32-1:0] FSM_fft_64_stage_1_0_t1132;
reg [6-1:0] FSM_fft_64_stage_1_0_t1133;
reg [32-1:0] FSM_fft_64_stage_1_0_t1134;
reg [33-1:0] FSM_fft_64_stage_1_0_t1135;
reg [32-1:0] FSM_fft_64_stage_1_0_t1136;
reg [2048-1:0] FSM_fft_64_stage_1_0_t1137;
reg [64-1:0] FSM_fft_64_stage_1_0_t1138;
reg [32-1:0] FSM_fft_64_stage_1_0_t1139;
reg [33-1:0] FSM_fft_64_stage_1_0_t1140;
reg [32-1:0] FSM_fft_64_stage_1_0_t1141;
reg [6-1:0] FSM_fft_64_stage_1_0_t1142;
reg [2048-1:0] FSM_fft_64_stage_1_0_t1143;
reg [64-1:0] FSM_fft_64_stage_1_0_t1144;
reg [32-1:0] FSM_fft_64_stage_1_0_t1145;
reg [6-1:0] FSM_fft_64_stage_1_0_t1146;
reg [64-1:0] FSM_fft_64_stage_1_0_t1147;
reg [32-1:0] FSM_fft_64_stage_1_0_t1148;
reg [6-1:0] FSM_fft_64_stage_1_0_t1149;
reg [32-1:0] FSM_fft_64_stage_1_0_t1150;
reg [64-1:0] FSM_fft_64_stage_1_0_t1151;
reg [32-1:0] FSM_fft_64_stage_1_0_t1152;
reg [33-1:0] FSM_fft_64_stage_1_0_t1153;
reg [32-1:0] FSM_fft_64_stage_1_0_t1154;
reg [6-1:0] FSM_fft_64_stage_1_0_t1155;
reg [32-1:0] FSM_fft_64_stage_1_0_t1156;
reg [33-1:0] FSM_fft_64_stage_1_0_t1157;
reg [32-1:0] FSM_fft_64_stage_1_0_t1158;
reg [2048-1:0] FSM_fft_64_stage_1_0_t1159;
reg [64-1:0] FSM_fft_64_stage_1_0_t1160;
reg [32-1:0] FSM_fft_64_stage_1_0_t1161;
reg [33-1:0] FSM_fft_64_stage_1_0_t1162;
reg [32-1:0] FSM_fft_64_stage_1_0_t1163;
reg [6-1:0] FSM_fft_64_stage_1_0_t1164;
reg [2048-1:0] FSM_fft_64_stage_1_0_t1165;
reg [64-1:0] FSM_fft_64_stage_1_0_t1166;
reg [32-1:0] FSM_fft_64_stage_1_0_t1167;
reg [6-1:0] FSM_fft_64_stage_1_0_t1168;
reg [64-1:0] FSM_fft_64_stage_1_0_t1169;
reg [32-1:0] FSM_fft_64_stage_1_0_t1170;
reg [6-1:0] FSM_fft_64_stage_1_0_t1171;
reg [32-1:0] FSM_fft_64_stage_1_0_t1172;
reg [64-1:0] FSM_fft_64_stage_1_0_t1173;
reg [32-1:0] FSM_fft_64_stage_1_0_t1174;
reg [33-1:0] FSM_fft_64_stage_1_0_t1175;
reg [32-1:0] FSM_fft_64_stage_1_0_t1176;
reg [6-1:0] FSM_fft_64_stage_1_0_t1177;
reg [32-1:0] FSM_fft_64_stage_1_0_t1178;
reg [33-1:0] FSM_fft_64_stage_1_0_t1179;
reg [32-1:0] FSM_fft_64_stage_1_0_t1180;
reg [2048-1:0] FSM_fft_64_stage_1_0_t1181;
reg [64-1:0] FSM_fft_64_stage_1_0_t1182;
reg [32-1:0] FSM_fft_64_stage_1_0_t1183;
reg [33-1:0] FSM_fft_64_stage_1_0_t1184;
reg [32-1:0] FSM_fft_64_stage_1_0_t1185;
reg [6-1:0] FSM_fft_64_stage_1_0_t1186;
reg [2048-1:0] FSM_fft_64_stage_1_0_t1187;
reg [64-1:0] FSM_fft_64_stage_1_0_t1188;
reg [32-1:0] FSM_fft_64_stage_1_0_t1189;
reg [6-1:0] FSM_fft_64_stage_1_0_t1190;
reg [64-1:0] FSM_fft_64_stage_1_0_t1191;
reg [32-1:0] FSM_fft_64_stage_1_0_t1192;
reg [6-1:0] FSM_fft_64_stage_1_0_t1193;
reg [32-1:0] FSM_fft_64_stage_1_0_t1194;
reg [64-1:0] FSM_fft_64_stage_1_0_t1195;
reg [32-1:0] FSM_fft_64_stage_1_0_t1196;
reg [33-1:0] FSM_fft_64_stage_1_0_t1197;
reg [32-1:0] FSM_fft_64_stage_1_0_t1198;
reg [6-1:0] FSM_fft_64_stage_1_0_t1199;
reg [32-1:0] FSM_fft_64_stage_1_0_t1200;
reg [33-1:0] FSM_fft_64_stage_1_0_t1201;
reg [32-1:0] FSM_fft_64_stage_1_0_t1202;
reg [2048-1:0] FSM_fft_64_stage_1_0_t1203;
reg [64-1:0] FSM_fft_64_stage_1_0_t1204;
reg [32-1:0] FSM_fft_64_stage_1_0_t1205;
reg [33-1:0] FSM_fft_64_stage_1_0_t1206;
reg [32-1:0] FSM_fft_64_stage_1_0_t1207;
reg [6-1:0] FSM_fft_64_stage_1_0_t1208;
reg [2048-1:0] FSM_fft_64_stage_1_0_t1209;
reg [64-1:0] FSM_fft_64_stage_1_0_t1210;
reg [32-1:0] FSM_fft_64_stage_1_0_t1211;
reg [6-1:0] FSM_fft_64_stage_1_0_t1212;
reg [64-1:0] FSM_fft_64_stage_1_0_t1213;
reg [32-1:0] FSM_fft_64_stage_1_0_t1214;
reg [6-1:0] FSM_fft_64_stage_1_0_t1215;
reg [32-1:0] FSM_fft_64_stage_1_0_t1216;
reg [64-1:0] FSM_fft_64_stage_1_0_t1217;
reg [32-1:0] FSM_fft_64_stage_1_0_t1218;
reg [33-1:0] FSM_fft_64_stage_1_0_t1219;
reg [32-1:0] FSM_fft_64_stage_1_0_t1220;
reg [6-1:0] FSM_fft_64_stage_1_0_t1221;
reg [32-1:0] FSM_fft_64_stage_1_0_t1222;
reg [33-1:0] FSM_fft_64_stage_1_0_t1223;
reg [32-1:0] FSM_fft_64_stage_1_0_t1224;
reg [2048-1:0] FSM_fft_64_stage_1_0_t1225;
reg [64-1:0] FSM_fft_64_stage_1_0_t1226;
reg [32-1:0] FSM_fft_64_stage_1_0_t1227;
reg [33-1:0] FSM_fft_64_stage_1_0_t1228;
reg [32-1:0] FSM_fft_64_stage_1_0_t1229;
reg [6-1:0] FSM_fft_64_stage_1_0_t1230;
reg [2048-1:0] FSM_fft_64_stage_1_0_t1231;
reg [64-1:0] FSM_fft_64_stage_1_0_t1232;
reg [32-1:0] FSM_fft_64_stage_1_0_t1233;
reg [6-1:0] FSM_fft_64_stage_1_0_t1234;
reg [64-1:0] FSM_fft_64_stage_1_0_t1235;
reg [32-1:0] FSM_fft_64_stage_1_0_t1236;
reg [6-1:0] FSM_fft_64_stage_1_0_t1237;
reg [32-1:0] FSM_fft_64_stage_1_0_t1238;
reg [64-1:0] FSM_fft_64_stage_1_0_t1239;
reg [32-1:0] FSM_fft_64_stage_1_0_t1240;
reg [33-1:0] FSM_fft_64_stage_1_0_t1241;
reg [32-1:0] FSM_fft_64_stage_1_0_t1242;
reg [6-1:0] FSM_fft_64_stage_1_0_t1243;
reg [32-1:0] FSM_fft_64_stage_1_0_t1244;
reg [33-1:0] FSM_fft_64_stage_1_0_t1245;
reg [32-1:0] FSM_fft_64_stage_1_0_t1246;
reg [2048-1:0] FSM_fft_64_stage_1_0_t1247;
reg [64-1:0] FSM_fft_64_stage_1_0_t1248;
reg [32-1:0] FSM_fft_64_stage_1_0_t1249;
reg [33-1:0] FSM_fft_64_stage_1_0_t1250;
reg [32-1:0] FSM_fft_64_stage_1_0_t1251;
reg [6-1:0] FSM_fft_64_stage_1_0_t1252;
reg [2048-1:0] FSM_fft_64_stage_1_0_t1253;
reg [64-1:0] FSM_fft_64_stage_1_0_t1254;
reg [32-1:0] FSM_fft_64_stage_1_0_t1255;
reg [6-1:0] FSM_fft_64_stage_1_0_t1256;
reg [64-1:0] FSM_fft_64_stage_1_0_t1257;
reg [32-1:0] FSM_fft_64_stage_1_0_t1258;
reg [6-1:0] FSM_fft_64_stage_1_0_t1259;
reg [32-1:0] FSM_fft_64_stage_1_0_t1260;
reg [64-1:0] FSM_fft_64_stage_1_0_t1261;
reg [32-1:0] FSM_fft_64_stage_1_0_t1262;
reg [33-1:0] FSM_fft_64_stage_1_0_t1263;
reg [32-1:0] FSM_fft_64_stage_1_0_t1264;
reg [6-1:0] FSM_fft_64_stage_1_0_t1265;
reg [32-1:0] FSM_fft_64_stage_1_0_t1266;
reg [33-1:0] FSM_fft_64_stage_1_0_t1267;
reg [32-1:0] FSM_fft_64_stage_1_0_t1268;
reg [2048-1:0] FSM_fft_64_stage_1_0_t1269;
reg [64-1:0] FSM_fft_64_stage_1_0_t1270;
reg [32-1:0] FSM_fft_64_stage_1_0_t1271;
reg [33-1:0] FSM_fft_64_stage_1_0_t1272;
reg [32-1:0] FSM_fft_64_stage_1_0_t1273;
reg [6-1:0] FSM_fft_64_stage_1_0_t1274;
reg [2048-1:0] FSM_fft_64_stage_1_0_t1275;
reg [64-1:0] FSM_fft_64_stage_1_0_t1276;
reg [32-1:0] FSM_fft_64_stage_1_0_t1277;
reg [6-1:0] FSM_fft_64_stage_1_0_t1278;
reg [64-1:0] FSM_fft_64_stage_1_0_t1279;
reg [32-1:0] FSM_fft_64_stage_1_0_t1280;
reg [6-1:0] FSM_fft_64_stage_1_0_t1281;
reg [32-1:0] FSM_fft_64_stage_1_0_t1282;
reg [64-1:0] FSM_fft_64_stage_1_0_t1283;
reg [32-1:0] FSM_fft_64_stage_1_0_t1284;
reg [33-1:0] FSM_fft_64_stage_1_0_t1285;
reg [32-1:0] FSM_fft_64_stage_1_0_t1286;
reg [6-1:0] FSM_fft_64_stage_1_0_t1287;
reg [32-1:0] FSM_fft_64_stage_1_0_t1288;
reg [33-1:0] FSM_fft_64_stage_1_0_t1289;
reg [32-1:0] FSM_fft_64_stage_1_0_t1290;
reg [2048-1:0] FSM_fft_64_stage_1_0_t1291;
reg [64-1:0] FSM_fft_64_stage_1_0_t1292;
reg [32-1:0] FSM_fft_64_stage_1_0_t1293;
reg [33-1:0] FSM_fft_64_stage_1_0_t1294;
reg [32-1:0] FSM_fft_64_stage_1_0_t1295;
reg [6-1:0] FSM_fft_64_stage_1_0_t1296;
reg [2048-1:0] FSM_fft_64_stage_1_0_t1297;
reg [64-1:0] FSM_fft_64_stage_1_0_t1298;
reg [32-1:0] FSM_fft_64_stage_1_0_t1299;
reg [6-1:0] FSM_fft_64_stage_1_0_t1300;
reg [64-1:0] FSM_fft_64_stage_1_0_t1301;
reg [32-1:0] FSM_fft_64_stage_1_0_t1302;
reg [6-1:0] FSM_fft_64_stage_1_0_t1303;
reg [32-1:0] FSM_fft_64_stage_1_0_t1304;
reg [64-1:0] FSM_fft_64_stage_1_0_t1305;
reg [32-1:0] FSM_fft_64_stage_1_0_t1306;
reg [33-1:0] FSM_fft_64_stage_1_0_t1307;
reg [32-1:0] FSM_fft_64_stage_1_0_t1308;
reg [6-1:0] FSM_fft_64_stage_1_0_t1309;
reg [32-1:0] FSM_fft_64_stage_1_0_t1310;
reg [33-1:0] FSM_fft_64_stage_1_0_t1311;
reg [32-1:0] FSM_fft_64_stage_1_0_t1312;
reg [2048-1:0] FSM_fft_64_stage_1_0_t1313;
reg [64-1:0] FSM_fft_64_stage_1_0_t1314;
reg [32-1:0] FSM_fft_64_stage_1_0_t1315;
reg [33-1:0] FSM_fft_64_stage_1_0_t1316;
reg [32-1:0] FSM_fft_64_stage_1_0_t1317;
reg [6-1:0] FSM_fft_64_stage_1_0_t1318;
reg [2048-1:0] FSM_fft_64_stage_1_0_t1319;
reg [64-1:0] FSM_fft_64_stage_1_0_t1320;
reg [32-1:0] FSM_fft_64_stage_1_0_t1321;
reg [6-1:0] FSM_fft_64_stage_1_0_t1322;
reg [64-1:0] FSM_fft_64_stage_1_0_t1323;
reg [32-1:0] FSM_fft_64_stage_1_0_t1324;
reg [6-1:0] FSM_fft_64_stage_1_0_t1325;
reg [32-1:0] FSM_fft_64_stage_1_0_t1326;
reg [64-1:0] FSM_fft_64_stage_1_0_t1327;
reg [32-1:0] FSM_fft_64_stage_1_0_t1328;
reg [33-1:0] FSM_fft_64_stage_1_0_t1329;
reg [32-1:0] FSM_fft_64_stage_1_0_t1330;
reg [6-1:0] FSM_fft_64_stage_1_0_t1331;
reg [32-1:0] FSM_fft_64_stage_1_0_t1332;
reg [33-1:0] FSM_fft_64_stage_1_0_t1333;
reg [32-1:0] FSM_fft_64_stage_1_0_t1334;
reg [2048-1:0] FSM_fft_64_stage_1_0_t1335;
reg [64-1:0] FSM_fft_64_stage_1_0_t1336;
reg [32-1:0] FSM_fft_64_stage_1_0_t1337;
reg [33-1:0] FSM_fft_64_stage_1_0_t1338;
reg [32-1:0] FSM_fft_64_stage_1_0_t1339;
reg [6-1:0] FSM_fft_64_stage_1_0_t1340;
reg [2048-1:0] FSM_fft_64_stage_1_0_t1341;
reg [64-1:0] FSM_fft_64_stage_1_0_t1342;
reg [32-1:0] FSM_fft_64_stage_1_0_t1343;
reg [6-1:0] FSM_fft_64_stage_1_0_t1344;
reg [64-1:0] FSM_fft_64_stage_1_0_t1345;
reg [32-1:0] FSM_fft_64_stage_1_0_t1346;
reg [6-1:0] FSM_fft_64_stage_1_0_t1347;
reg [32-1:0] FSM_fft_64_stage_1_0_t1348;
reg [64-1:0] FSM_fft_64_stage_1_0_t1349;
reg [32-1:0] FSM_fft_64_stage_1_0_t1350;
reg [33-1:0] FSM_fft_64_stage_1_0_t1351;
reg [32-1:0] FSM_fft_64_stage_1_0_t1352;
reg [6-1:0] FSM_fft_64_stage_1_0_t1353;
reg [32-1:0] FSM_fft_64_stage_1_0_t1354;
reg [33-1:0] FSM_fft_64_stage_1_0_t1355;
reg [32-1:0] FSM_fft_64_stage_1_0_t1356;
reg [2048-1:0] FSM_fft_64_stage_1_0_t1357;
reg [64-1:0] FSM_fft_64_stage_1_0_t1358;
reg [32-1:0] FSM_fft_64_stage_1_0_t1359;
reg [33-1:0] FSM_fft_64_stage_1_0_t1360;
reg [32-1:0] FSM_fft_64_stage_1_0_t1361;
reg [6-1:0] FSM_fft_64_stage_1_0_t1362;
reg [2048-1:0] FSM_fft_64_stage_1_0_t1363;
reg [64-1:0] FSM_fft_64_stage_1_0_t1364;
reg [32-1:0] FSM_fft_64_stage_1_0_t1365;
reg [6-1:0] FSM_fft_64_stage_1_0_t1366;
reg [64-1:0] FSM_fft_64_stage_1_0_t1367;
reg [32-1:0] FSM_fft_64_stage_1_0_t1368;
reg [6-1:0] FSM_fft_64_stage_1_0_t1369;
reg [32-1:0] FSM_fft_64_stage_1_0_t1370;
reg [64-1:0] FSM_fft_64_stage_1_0_t1371;
reg [32-1:0] FSM_fft_64_stage_1_0_t1372;
reg [33-1:0] FSM_fft_64_stage_1_0_t1373;
reg [32-1:0] FSM_fft_64_stage_1_0_t1374;
reg [6-1:0] FSM_fft_64_stage_1_0_t1375;
reg [32-1:0] FSM_fft_64_stage_1_0_t1376;
reg [33-1:0] FSM_fft_64_stage_1_0_t1377;
reg [32-1:0] FSM_fft_64_stage_1_0_t1378;
reg [2048-1:0] FSM_fft_64_stage_1_0_t1379;
reg [64-1:0] FSM_fft_64_stage_1_0_t1380;
reg [32-1:0] FSM_fft_64_stage_1_0_t1381;
reg [33-1:0] FSM_fft_64_stage_1_0_t1382;
reg [32-1:0] FSM_fft_64_stage_1_0_t1383;
reg [6-1:0] FSM_fft_64_stage_1_0_t1384;
reg [2048-1:0] FSM_fft_64_stage_1_0_t1385;
reg [64-1:0] FSM_fft_64_stage_1_0_t1386;
reg [32-1:0] FSM_fft_64_stage_1_0_t1387;
reg [6-1:0] FSM_fft_64_stage_1_0_t1388;
reg [64-1:0] FSM_fft_64_stage_1_0_t1389;
reg [32-1:0] FSM_fft_64_stage_1_0_t1390;
reg [6-1:0] FSM_fft_64_stage_1_0_t1391;
reg [32-1:0] FSM_fft_64_stage_1_0_t1392;
reg [64-1:0] FSM_fft_64_stage_1_0_t1393;
reg [32-1:0] FSM_fft_64_stage_1_0_t1394;
reg [33-1:0] FSM_fft_64_stage_1_0_t1395;
reg [32-1:0] FSM_fft_64_stage_1_0_t1396;
reg [6-1:0] FSM_fft_64_stage_1_0_t1397;
reg [32-1:0] FSM_fft_64_stage_1_0_t1398;
reg [33-1:0] FSM_fft_64_stage_1_0_t1399;
reg [32-1:0] FSM_fft_64_stage_1_0_t1400;
reg [2048-1:0] FSM_fft_64_stage_1_0_t1401;
reg [64-1:0] FSM_fft_64_stage_1_0_t1402;
reg [32-1:0] FSM_fft_64_stage_1_0_t1403;
reg [33-1:0] FSM_fft_64_stage_1_0_t1404;
reg [32-1:0] FSM_fft_64_stage_1_0_t1405;
reg [6-1:0] FSM_fft_64_stage_1_0_t1406;
reg [2048-1:0] FSM_fft_64_stage_1_0_t1407;

assign FSM_fft_64_stage_1_0_out_valid = 1'b1;
/*
    Wiring by fft_64_stage_1
*/
assign i_ready = FSM_fft_64_stage_1_0_in_ready;
assign o_data_out_real = FSM_fft_64_stage_1_0_t703;
assign o_data_out_imag = FSM_fft_64_stage_1_0_t1407;
assign o_valid = FSM_fft_64_stage_1_0_out_valid;
/* End wiring by fft_64_stage_1 */


initial begin
    FSM_fft_64_stage_1_0_t0 = 32'b00000000000000000000000000000010 * 32'b0;
    FSM_fft_64_stage_1_0_t1 = FSM_fft_64_stage_1_0_t0[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t2 = FSM_fft_64_stage_1_0_t1[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t3 = 32'b00000000000000000000000000000010 * 32'b0;
    FSM_fft_64_stage_1_0_t4 = FSM_fft_64_stage_1_0_t3[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t5 = FSM_fft_64_stage_1_0_t4[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t6 = i_data_in_real[FSM_fft_64_stage_1_0_t5 * 32 +: 32];
    FSM_fft_64_stage_1_0_t7 = 32'b00000000000000000000000000000010 * 32'b0;
    FSM_fft_64_stage_1_0_t8 = FSM_fft_64_stage_1_0_t7[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t9 = FSM_fft_64_stage_1_0_t8 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t10 = FSM_fft_64_stage_1_0_t9[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t11 = FSM_fft_64_stage_1_0_t10[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t12 = i_data_in_real[FSM_fft_64_stage_1_0_t11 * 32 +: 32];
    FSM_fft_64_stage_1_0_t13 = FSM_fft_64_stage_1_0_t6 + FSM_fft_64_stage_1_0_t12;
    FSM_fft_64_stage_1_0_t14 = FSM_fft_64_stage_1_0_t13[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t15 = 2048'b0;
    FSM_fft_64_stage_1_0_t15[FSM_fft_64_stage_1_0_t2 * 32 +: 32] = FSM_fft_64_stage_1_0_t14;
    FSM_fft_64_stage_1_0_t16 = 32'b00000000000000000000000000000010 * 32'b0;
    FSM_fft_64_stage_1_0_t17 = FSM_fft_64_stage_1_0_t16[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t18 = FSM_fft_64_stage_1_0_t17 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t19 = FSM_fft_64_stage_1_0_t18[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t20 = FSM_fft_64_stage_1_0_t19[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t21 = FSM_fft_64_stage_1_0_t15;
    FSM_fft_64_stage_1_0_t21[FSM_fft_64_stage_1_0_t20 * 32 +: 32] = FSM_fft_64_stage_1_0_t6 - FSM_fft_64_stage_1_0_t12;
    FSM_fft_64_stage_1_0_t22 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t23 = FSM_fft_64_stage_1_0_t22[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t24 = FSM_fft_64_stage_1_0_t23[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t25 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t26 = FSM_fft_64_stage_1_0_t25[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t27 = FSM_fft_64_stage_1_0_t26[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t28 = i_data_in_real[FSM_fft_64_stage_1_0_t27 * 32 +: 32];
    FSM_fft_64_stage_1_0_t29 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t30 = FSM_fft_64_stage_1_0_t29[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t31 = FSM_fft_64_stage_1_0_t30 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t32 = FSM_fft_64_stage_1_0_t31[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t33 = FSM_fft_64_stage_1_0_t32[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t34 = i_data_in_real[FSM_fft_64_stage_1_0_t33 * 32 +: 32];
    FSM_fft_64_stage_1_0_t35 = FSM_fft_64_stage_1_0_t28 + FSM_fft_64_stage_1_0_t34;
    FSM_fft_64_stage_1_0_t36 = FSM_fft_64_stage_1_0_t35[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t37 = FSM_fft_64_stage_1_0_t21;
    FSM_fft_64_stage_1_0_t37[FSM_fft_64_stage_1_0_t24 * 32 +: 32] = FSM_fft_64_stage_1_0_t36;
    FSM_fft_64_stage_1_0_t38 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t39 = FSM_fft_64_stage_1_0_t38[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t40 = FSM_fft_64_stage_1_0_t39 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t41 = FSM_fft_64_stage_1_0_t40[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t42 = FSM_fft_64_stage_1_0_t41[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t43 = FSM_fft_64_stage_1_0_t37;
    FSM_fft_64_stage_1_0_t43[FSM_fft_64_stage_1_0_t42 * 32 +: 32] = FSM_fft_64_stage_1_0_t28 - FSM_fft_64_stage_1_0_t34;
    FSM_fft_64_stage_1_0_t44 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_1_0_t45 = FSM_fft_64_stage_1_0_t44[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t46 = FSM_fft_64_stage_1_0_t45[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t47 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_1_0_t48 = FSM_fft_64_stage_1_0_t47[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t49 = FSM_fft_64_stage_1_0_t48[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t50 = i_data_in_real[FSM_fft_64_stage_1_0_t49 * 32 +: 32];
    FSM_fft_64_stage_1_0_t51 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_1_0_t52 = FSM_fft_64_stage_1_0_t51[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t53 = FSM_fft_64_stage_1_0_t52 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t54 = FSM_fft_64_stage_1_0_t53[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t55 = FSM_fft_64_stage_1_0_t54[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t56 = i_data_in_real[FSM_fft_64_stage_1_0_t55 * 32 +: 32];
    FSM_fft_64_stage_1_0_t57 = FSM_fft_64_stage_1_0_t50 + FSM_fft_64_stage_1_0_t56;
    FSM_fft_64_stage_1_0_t58 = FSM_fft_64_stage_1_0_t57[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t59 = FSM_fft_64_stage_1_0_t43;
    FSM_fft_64_stage_1_0_t59[FSM_fft_64_stage_1_0_t46 * 32 +: 32] = FSM_fft_64_stage_1_0_t58;
    FSM_fft_64_stage_1_0_t60 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_1_0_t61 = FSM_fft_64_stage_1_0_t60[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t62 = FSM_fft_64_stage_1_0_t61 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t63 = FSM_fft_64_stage_1_0_t62[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t64 = FSM_fft_64_stage_1_0_t63[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t65 = FSM_fft_64_stage_1_0_t59;
    FSM_fft_64_stage_1_0_t65[FSM_fft_64_stage_1_0_t64 * 32 +: 32] = FSM_fft_64_stage_1_0_t50 - FSM_fft_64_stage_1_0_t56;
    FSM_fft_64_stage_1_0_t66 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_1_0_t67 = FSM_fft_64_stage_1_0_t66[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t68 = FSM_fft_64_stage_1_0_t67[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t69 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_1_0_t70 = FSM_fft_64_stage_1_0_t69[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t71 = FSM_fft_64_stage_1_0_t70[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t72 = i_data_in_real[FSM_fft_64_stage_1_0_t71 * 32 +: 32];
    FSM_fft_64_stage_1_0_t73 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_1_0_t74 = FSM_fft_64_stage_1_0_t73[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t75 = FSM_fft_64_stage_1_0_t74 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t76 = FSM_fft_64_stage_1_0_t75[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t77 = FSM_fft_64_stage_1_0_t76[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t78 = i_data_in_real[FSM_fft_64_stage_1_0_t77 * 32 +: 32];
    FSM_fft_64_stage_1_0_t79 = FSM_fft_64_stage_1_0_t72 + FSM_fft_64_stage_1_0_t78;
    FSM_fft_64_stage_1_0_t80 = FSM_fft_64_stage_1_0_t79[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t81 = FSM_fft_64_stage_1_0_t65;
    FSM_fft_64_stage_1_0_t81[FSM_fft_64_stage_1_0_t68 * 32 +: 32] = FSM_fft_64_stage_1_0_t80;
    FSM_fft_64_stage_1_0_t82 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_1_0_t83 = FSM_fft_64_stage_1_0_t82[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t84 = FSM_fft_64_stage_1_0_t83 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t85 = FSM_fft_64_stage_1_0_t84[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t86 = FSM_fft_64_stage_1_0_t85[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t87 = FSM_fft_64_stage_1_0_t81;
    FSM_fft_64_stage_1_0_t87[FSM_fft_64_stage_1_0_t86 * 32 +: 32] = FSM_fft_64_stage_1_0_t72 - FSM_fft_64_stage_1_0_t78;
    FSM_fft_64_stage_1_0_t88 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000100;
    FSM_fft_64_stage_1_0_t89 = FSM_fft_64_stage_1_0_t88[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t90 = FSM_fft_64_stage_1_0_t89[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t91 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000100;
    FSM_fft_64_stage_1_0_t92 = FSM_fft_64_stage_1_0_t91[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t93 = FSM_fft_64_stage_1_0_t92[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t94 = i_data_in_real[FSM_fft_64_stage_1_0_t93 * 32 +: 32];
    FSM_fft_64_stage_1_0_t95 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000100;
    FSM_fft_64_stage_1_0_t96 = FSM_fft_64_stage_1_0_t95[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t97 = FSM_fft_64_stage_1_0_t96 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t98 = FSM_fft_64_stage_1_0_t97[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t99 = FSM_fft_64_stage_1_0_t98[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t100 = i_data_in_real[FSM_fft_64_stage_1_0_t99 * 32 +: 32];
    FSM_fft_64_stage_1_0_t101 = FSM_fft_64_stage_1_0_t94 + FSM_fft_64_stage_1_0_t100;
    FSM_fft_64_stage_1_0_t102 = FSM_fft_64_stage_1_0_t101[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t103 = FSM_fft_64_stage_1_0_t87;
    FSM_fft_64_stage_1_0_t103[FSM_fft_64_stage_1_0_t90 * 32 +: 32] = FSM_fft_64_stage_1_0_t102;
    FSM_fft_64_stage_1_0_t104 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000100;
    FSM_fft_64_stage_1_0_t105 = FSM_fft_64_stage_1_0_t104[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t106 = FSM_fft_64_stage_1_0_t105 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t107 = FSM_fft_64_stage_1_0_t106[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t108 = FSM_fft_64_stage_1_0_t107[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t109 = FSM_fft_64_stage_1_0_t103;
    FSM_fft_64_stage_1_0_t109[FSM_fft_64_stage_1_0_t108 * 32 +: 32] = FSM_fft_64_stage_1_0_t94 - FSM_fft_64_stage_1_0_t100;
    FSM_fft_64_stage_1_0_t110 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000101;
    FSM_fft_64_stage_1_0_t111 = FSM_fft_64_stage_1_0_t110[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t112 = FSM_fft_64_stage_1_0_t111[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t113 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000101;
    FSM_fft_64_stage_1_0_t114 = FSM_fft_64_stage_1_0_t113[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t115 = FSM_fft_64_stage_1_0_t114[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t116 = i_data_in_real[FSM_fft_64_stage_1_0_t115 * 32 +: 32];
    FSM_fft_64_stage_1_0_t117 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000101;
    FSM_fft_64_stage_1_0_t118 = FSM_fft_64_stage_1_0_t117[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t119 = FSM_fft_64_stage_1_0_t118 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t120 = FSM_fft_64_stage_1_0_t119[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t121 = FSM_fft_64_stage_1_0_t120[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t122 = i_data_in_real[FSM_fft_64_stage_1_0_t121 * 32 +: 32];
    FSM_fft_64_stage_1_0_t123 = FSM_fft_64_stage_1_0_t116 + FSM_fft_64_stage_1_0_t122;
    FSM_fft_64_stage_1_0_t124 = FSM_fft_64_stage_1_0_t123[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t125 = FSM_fft_64_stage_1_0_t109;
    FSM_fft_64_stage_1_0_t125[FSM_fft_64_stage_1_0_t112 * 32 +: 32] = FSM_fft_64_stage_1_0_t124;
    FSM_fft_64_stage_1_0_t126 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000101;
    FSM_fft_64_stage_1_0_t127 = FSM_fft_64_stage_1_0_t126[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t128 = FSM_fft_64_stage_1_0_t127 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t129 = FSM_fft_64_stage_1_0_t128[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t130 = FSM_fft_64_stage_1_0_t129[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t131 = FSM_fft_64_stage_1_0_t125;
    FSM_fft_64_stage_1_0_t131[FSM_fft_64_stage_1_0_t130 * 32 +: 32] = FSM_fft_64_stage_1_0_t116 - FSM_fft_64_stage_1_0_t122;
    FSM_fft_64_stage_1_0_t132 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000110;
    FSM_fft_64_stage_1_0_t133 = FSM_fft_64_stage_1_0_t132[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t134 = FSM_fft_64_stage_1_0_t133[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t135 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000110;
    FSM_fft_64_stage_1_0_t136 = FSM_fft_64_stage_1_0_t135[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t137 = FSM_fft_64_stage_1_0_t136[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t138 = i_data_in_real[FSM_fft_64_stage_1_0_t137 * 32 +: 32];
    FSM_fft_64_stage_1_0_t139 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000110;
    FSM_fft_64_stage_1_0_t140 = FSM_fft_64_stage_1_0_t139[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t141 = FSM_fft_64_stage_1_0_t140 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t142 = FSM_fft_64_stage_1_0_t141[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t143 = FSM_fft_64_stage_1_0_t142[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t144 = i_data_in_real[FSM_fft_64_stage_1_0_t143 * 32 +: 32];
    FSM_fft_64_stage_1_0_t145 = FSM_fft_64_stage_1_0_t138 + FSM_fft_64_stage_1_0_t144;
    FSM_fft_64_stage_1_0_t146 = FSM_fft_64_stage_1_0_t145[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t147 = FSM_fft_64_stage_1_0_t131;
    FSM_fft_64_stage_1_0_t147[FSM_fft_64_stage_1_0_t134 * 32 +: 32] = FSM_fft_64_stage_1_0_t146;
    FSM_fft_64_stage_1_0_t148 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000110;
    FSM_fft_64_stage_1_0_t149 = FSM_fft_64_stage_1_0_t148[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t150 = FSM_fft_64_stage_1_0_t149 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t151 = FSM_fft_64_stage_1_0_t150[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t152 = FSM_fft_64_stage_1_0_t151[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t153 = FSM_fft_64_stage_1_0_t147;
    FSM_fft_64_stage_1_0_t153[FSM_fft_64_stage_1_0_t152 * 32 +: 32] = FSM_fft_64_stage_1_0_t138 - FSM_fft_64_stage_1_0_t144;
    FSM_fft_64_stage_1_0_t154 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000111;
    FSM_fft_64_stage_1_0_t155 = FSM_fft_64_stage_1_0_t154[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t156 = FSM_fft_64_stage_1_0_t155[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t157 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000111;
    FSM_fft_64_stage_1_0_t158 = FSM_fft_64_stage_1_0_t157[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t159 = FSM_fft_64_stage_1_0_t158[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t160 = i_data_in_real[FSM_fft_64_stage_1_0_t159 * 32 +: 32];
    FSM_fft_64_stage_1_0_t161 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000111;
    FSM_fft_64_stage_1_0_t162 = FSM_fft_64_stage_1_0_t161[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t163 = FSM_fft_64_stage_1_0_t162 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t164 = FSM_fft_64_stage_1_0_t163[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t165 = FSM_fft_64_stage_1_0_t164[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t166 = i_data_in_real[FSM_fft_64_stage_1_0_t165 * 32 +: 32];
    FSM_fft_64_stage_1_0_t167 = FSM_fft_64_stage_1_0_t160 + FSM_fft_64_stage_1_0_t166;
    FSM_fft_64_stage_1_0_t168 = FSM_fft_64_stage_1_0_t167[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t169 = FSM_fft_64_stage_1_0_t153;
    FSM_fft_64_stage_1_0_t169[FSM_fft_64_stage_1_0_t156 * 32 +: 32] = FSM_fft_64_stage_1_0_t168;
    FSM_fft_64_stage_1_0_t170 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000111;
    FSM_fft_64_stage_1_0_t171 = FSM_fft_64_stage_1_0_t170[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t172 = FSM_fft_64_stage_1_0_t171 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t173 = FSM_fft_64_stage_1_0_t172[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t174 = FSM_fft_64_stage_1_0_t173[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t175 = FSM_fft_64_stage_1_0_t169;
    FSM_fft_64_stage_1_0_t175[FSM_fft_64_stage_1_0_t174 * 32 +: 32] = FSM_fft_64_stage_1_0_t160 - FSM_fft_64_stage_1_0_t166;
    FSM_fft_64_stage_1_0_t176 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001000;
    FSM_fft_64_stage_1_0_t177 = FSM_fft_64_stage_1_0_t176[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t178 = FSM_fft_64_stage_1_0_t177[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t179 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001000;
    FSM_fft_64_stage_1_0_t180 = FSM_fft_64_stage_1_0_t179[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t181 = FSM_fft_64_stage_1_0_t180[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t182 = i_data_in_real[FSM_fft_64_stage_1_0_t181 * 32 +: 32];
    FSM_fft_64_stage_1_0_t183 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001000;
    FSM_fft_64_stage_1_0_t184 = FSM_fft_64_stage_1_0_t183[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t185 = FSM_fft_64_stage_1_0_t184 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t186 = FSM_fft_64_stage_1_0_t185[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t187 = FSM_fft_64_stage_1_0_t186[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t188 = i_data_in_real[FSM_fft_64_stage_1_0_t187 * 32 +: 32];
    FSM_fft_64_stage_1_0_t189 = FSM_fft_64_stage_1_0_t182 + FSM_fft_64_stage_1_0_t188;
    FSM_fft_64_stage_1_0_t190 = FSM_fft_64_stage_1_0_t189[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t191 = FSM_fft_64_stage_1_0_t175;
    FSM_fft_64_stage_1_0_t191[FSM_fft_64_stage_1_0_t178 * 32 +: 32] = FSM_fft_64_stage_1_0_t190;
    FSM_fft_64_stage_1_0_t192 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001000;
    FSM_fft_64_stage_1_0_t193 = FSM_fft_64_stage_1_0_t192[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t194 = FSM_fft_64_stage_1_0_t193 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t195 = FSM_fft_64_stage_1_0_t194[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t196 = FSM_fft_64_stage_1_0_t195[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t197 = FSM_fft_64_stage_1_0_t191;
    FSM_fft_64_stage_1_0_t197[FSM_fft_64_stage_1_0_t196 * 32 +: 32] = FSM_fft_64_stage_1_0_t182 - FSM_fft_64_stage_1_0_t188;
    FSM_fft_64_stage_1_0_t198 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001001;
    FSM_fft_64_stage_1_0_t199 = FSM_fft_64_stage_1_0_t198[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t200 = FSM_fft_64_stage_1_0_t199[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t201 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001001;
    FSM_fft_64_stage_1_0_t202 = FSM_fft_64_stage_1_0_t201[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t203 = FSM_fft_64_stage_1_0_t202[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t204 = i_data_in_real[FSM_fft_64_stage_1_0_t203 * 32 +: 32];
    FSM_fft_64_stage_1_0_t205 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001001;
    FSM_fft_64_stage_1_0_t206 = FSM_fft_64_stage_1_0_t205[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t207 = FSM_fft_64_stage_1_0_t206 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t208 = FSM_fft_64_stage_1_0_t207[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t209 = FSM_fft_64_stage_1_0_t208[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t210 = i_data_in_real[FSM_fft_64_stage_1_0_t209 * 32 +: 32];
    FSM_fft_64_stage_1_0_t211 = FSM_fft_64_stage_1_0_t204 + FSM_fft_64_stage_1_0_t210;
    FSM_fft_64_stage_1_0_t212 = FSM_fft_64_stage_1_0_t211[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t213 = FSM_fft_64_stage_1_0_t197;
    FSM_fft_64_stage_1_0_t213[FSM_fft_64_stage_1_0_t200 * 32 +: 32] = FSM_fft_64_stage_1_0_t212;
    FSM_fft_64_stage_1_0_t214 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001001;
    FSM_fft_64_stage_1_0_t215 = FSM_fft_64_stage_1_0_t214[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t216 = FSM_fft_64_stage_1_0_t215 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t217 = FSM_fft_64_stage_1_0_t216[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t218 = FSM_fft_64_stage_1_0_t217[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t219 = FSM_fft_64_stage_1_0_t213;
    FSM_fft_64_stage_1_0_t219[FSM_fft_64_stage_1_0_t218 * 32 +: 32] = FSM_fft_64_stage_1_0_t204 - FSM_fft_64_stage_1_0_t210;
    FSM_fft_64_stage_1_0_t220 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001010;
    FSM_fft_64_stage_1_0_t221 = FSM_fft_64_stage_1_0_t220[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t222 = FSM_fft_64_stage_1_0_t221[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t223 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001010;
    FSM_fft_64_stage_1_0_t224 = FSM_fft_64_stage_1_0_t223[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t225 = FSM_fft_64_stage_1_0_t224[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t226 = i_data_in_real[FSM_fft_64_stage_1_0_t225 * 32 +: 32];
    FSM_fft_64_stage_1_0_t227 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001010;
    FSM_fft_64_stage_1_0_t228 = FSM_fft_64_stage_1_0_t227[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t229 = FSM_fft_64_stage_1_0_t228 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t230 = FSM_fft_64_stage_1_0_t229[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t231 = FSM_fft_64_stage_1_0_t230[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t232 = i_data_in_real[FSM_fft_64_stage_1_0_t231 * 32 +: 32];
    FSM_fft_64_stage_1_0_t233 = FSM_fft_64_stage_1_0_t226 + FSM_fft_64_stage_1_0_t232;
    FSM_fft_64_stage_1_0_t234 = FSM_fft_64_stage_1_0_t233[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t235 = FSM_fft_64_stage_1_0_t219;
    FSM_fft_64_stage_1_0_t235[FSM_fft_64_stage_1_0_t222 * 32 +: 32] = FSM_fft_64_stage_1_0_t234;
    FSM_fft_64_stage_1_0_t236 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001010;
    FSM_fft_64_stage_1_0_t237 = FSM_fft_64_stage_1_0_t236[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t238 = FSM_fft_64_stage_1_0_t237 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t239 = FSM_fft_64_stage_1_0_t238[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t240 = FSM_fft_64_stage_1_0_t239[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t241 = FSM_fft_64_stage_1_0_t235;
    FSM_fft_64_stage_1_0_t241[FSM_fft_64_stage_1_0_t240 * 32 +: 32] = FSM_fft_64_stage_1_0_t226 - FSM_fft_64_stage_1_0_t232;
    FSM_fft_64_stage_1_0_t242 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001011;
    FSM_fft_64_stage_1_0_t243 = FSM_fft_64_stage_1_0_t242[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t244 = FSM_fft_64_stage_1_0_t243[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t245 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001011;
    FSM_fft_64_stage_1_0_t246 = FSM_fft_64_stage_1_0_t245[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t247 = FSM_fft_64_stage_1_0_t246[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t248 = i_data_in_real[FSM_fft_64_stage_1_0_t247 * 32 +: 32];
    FSM_fft_64_stage_1_0_t249 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001011;
    FSM_fft_64_stage_1_0_t250 = FSM_fft_64_stage_1_0_t249[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t251 = FSM_fft_64_stage_1_0_t250 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t252 = FSM_fft_64_stage_1_0_t251[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t253 = FSM_fft_64_stage_1_0_t252[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t254 = i_data_in_real[FSM_fft_64_stage_1_0_t253 * 32 +: 32];
    FSM_fft_64_stage_1_0_t255 = FSM_fft_64_stage_1_0_t248 + FSM_fft_64_stage_1_0_t254;
    FSM_fft_64_stage_1_0_t256 = FSM_fft_64_stage_1_0_t255[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t257 = FSM_fft_64_stage_1_0_t241;
    FSM_fft_64_stage_1_0_t257[FSM_fft_64_stage_1_0_t244 * 32 +: 32] = FSM_fft_64_stage_1_0_t256;
    FSM_fft_64_stage_1_0_t258 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001011;
    FSM_fft_64_stage_1_0_t259 = FSM_fft_64_stage_1_0_t258[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t260 = FSM_fft_64_stage_1_0_t259 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t261 = FSM_fft_64_stage_1_0_t260[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t262 = FSM_fft_64_stage_1_0_t261[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t263 = FSM_fft_64_stage_1_0_t257;
    FSM_fft_64_stage_1_0_t263[FSM_fft_64_stage_1_0_t262 * 32 +: 32] = FSM_fft_64_stage_1_0_t248 - FSM_fft_64_stage_1_0_t254;
    FSM_fft_64_stage_1_0_t264 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001100;
    FSM_fft_64_stage_1_0_t265 = FSM_fft_64_stage_1_0_t264[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t266 = FSM_fft_64_stage_1_0_t265[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t267 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001100;
    FSM_fft_64_stage_1_0_t268 = FSM_fft_64_stage_1_0_t267[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t269 = FSM_fft_64_stage_1_0_t268[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t270 = i_data_in_real[FSM_fft_64_stage_1_0_t269 * 32 +: 32];
    FSM_fft_64_stage_1_0_t271 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001100;
    FSM_fft_64_stage_1_0_t272 = FSM_fft_64_stage_1_0_t271[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t273 = FSM_fft_64_stage_1_0_t272 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t274 = FSM_fft_64_stage_1_0_t273[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t275 = FSM_fft_64_stage_1_0_t274[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t276 = i_data_in_real[FSM_fft_64_stage_1_0_t275 * 32 +: 32];
    FSM_fft_64_stage_1_0_t277 = FSM_fft_64_stage_1_0_t270 + FSM_fft_64_stage_1_0_t276;
    FSM_fft_64_stage_1_0_t278 = FSM_fft_64_stage_1_0_t277[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t279 = FSM_fft_64_stage_1_0_t263;
    FSM_fft_64_stage_1_0_t279[FSM_fft_64_stage_1_0_t266 * 32 +: 32] = FSM_fft_64_stage_1_0_t278;
    FSM_fft_64_stage_1_0_t280 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001100;
    FSM_fft_64_stage_1_0_t281 = FSM_fft_64_stage_1_0_t280[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t282 = FSM_fft_64_stage_1_0_t281 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t283 = FSM_fft_64_stage_1_0_t282[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t284 = FSM_fft_64_stage_1_0_t283[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t285 = FSM_fft_64_stage_1_0_t279;
    FSM_fft_64_stage_1_0_t285[FSM_fft_64_stage_1_0_t284 * 32 +: 32] = FSM_fft_64_stage_1_0_t270 - FSM_fft_64_stage_1_0_t276;
    FSM_fft_64_stage_1_0_t286 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001101;
    FSM_fft_64_stage_1_0_t287 = FSM_fft_64_stage_1_0_t286[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t288 = FSM_fft_64_stage_1_0_t287[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t289 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001101;
    FSM_fft_64_stage_1_0_t290 = FSM_fft_64_stage_1_0_t289[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t291 = FSM_fft_64_stage_1_0_t290[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t292 = i_data_in_real[FSM_fft_64_stage_1_0_t291 * 32 +: 32];
    FSM_fft_64_stage_1_0_t293 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001101;
    FSM_fft_64_stage_1_0_t294 = FSM_fft_64_stage_1_0_t293[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t295 = FSM_fft_64_stage_1_0_t294 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t296 = FSM_fft_64_stage_1_0_t295[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t297 = FSM_fft_64_stage_1_0_t296[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t298 = i_data_in_real[FSM_fft_64_stage_1_0_t297 * 32 +: 32];
    FSM_fft_64_stage_1_0_t299 = FSM_fft_64_stage_1_0_t292 + FSM_fft_64_stage_1_0_t298;
    FSM_fft_64_stage_1_0_t300 = FSM_fft_64_stage_1_0_t299[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t301 = FSM_fft_64_stage_1_0_t285;
    FSM_fft_64_stage_1_0_t301[FSM_fft_64_stage_1_0_t288 * 32 +: 32] = FSM_fft_64_stage_1_0_t300;
    FSM_fft_64_stage_1_0_t302 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001101;
    FSM_fft_64_stage_1_0_t303 = FSM_fft_64_stage_1_0_t302[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t304 = FSM_fft_64_stage_1_0_t303 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t305 = FSM_fft_64_stage_1_0_t304[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t306 = FSM_fft_64_stage_1_0_t305[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t307 = FSM_fft_64_stage_1_0_t301;
    FSM_fft_64_stage_1_0_t307[FSM_fft_64_stage_1_0_t306 * 32 +: 32] = FSM_fft_64_stage_1_0_t292 - FSM_fft_64_stage_1_0_t298;
    FSM_fft_64_stage_1_0_t308 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001110;
    FSM_fft_64_stage_1_0_t309 = FSM_fft_64_stage_1_0_t308[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t310 = FSM_fft_64_stage_1_0_t309[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t311 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001110;
    FSM_fft_64_stage_1_0_t312 = FSM_fft_64_stage_1_0_t311[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t313 = FSM_fft_64_stage_1_0_t312[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t314 = i_data_in_real[FSM_fft_64_stage_1_0_t313 * 32 +: 32];
    FSM_fft_64_stage_1_0_t315 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001110;
    FSM_fft_64_stage_1_0_t316 = FSM_fft_64_stage_1_0_t315[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t317 = FSM_fft_64_stage_1_0_t316 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t318 = FSM_fft_64_stage_1_0_t317[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t319 = FSM_fft_64_stage_1_0_t318[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t320 = i_data_in_real[FSM_fft_64_stage_1_0_t319 * 32 +: 32];
    FSM_fft_64_stage_1_0_t321 = FSM_fft_64_stage_1_0_t314 + FSM_fft_64_stage_1_0_t320;
    FSM_fft_64_stage_1_0_t322 = FSM_fft_64_stage_1_0_t321[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t323 = FSM_fft_64_stage_1_0_t307;
    FSM_fft_64_stage_1_0_t323[FSM_fft_64_stage_1_0_t310 * 32 +: 32] = FSM_fft_64_stage_1_0_t322;
    FSM_fft_64_stage_1_0_t324 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001110;
    FSM_fft_64_stage_1_0_t325 = FSM_fft_64_stage_1_0_t324[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t326 = FSM_fft_64_stage_1_0_t325 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t327 = FSM_fft_64_stage_1_0_t326[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t328 = FSM_fft_64_stage_1_0_t327[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t329 = FSM_fft_64_stage_1_0_t323;
    FSM_fft_64_stage_1_0_t329[FSM_fft_64_stage_1_0_t328 * 32 +: 32] = FSM_fft_64_stage_1_0_t314 - FSM_fft_64_stage_1_0_t320;
    FSM_fft_64_stage_1_0_t330 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001111;
    FSM_fft_64_stage_1_0_t331 = FSM_fft_64_stage_1_0_t330[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t332 = FSM_fft_64_stage_1_0_t331[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t333 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001111;
    FSM_fft_64_stage_1_0_t334 = FSM_fft_64_stage_1_0_t333[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t335 = FSM_fft_64_stage_1_0_t334[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t336 = i_data_in_real[FSM_fft_64_stage_1_0_t335 * 32 +: 32];
    FSM_fft_64_stage_1_0_t337 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001111;
    FSM_fft_64_stage_1_0_t338 = FSM_fft_64_stage_1_0_t337[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t339 = FSM_fft_64_stage_1_0_t338 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t340 = FSM_fft_64_stage_1_0_t339[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t341 = FSM_fft_64_stage_1_0_t340[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t342 = i_data_in_real[FSM_fft_64_stage_1_0_t341 * 32 +: 32];
    FSM_fft_64_stage_1_0_t343 = FSM_fft_64_stage_1_0_t336 + FSM_fft_64_stage_1_0_t342;
    FSM_fft_64_stage_1_0_t344 = FSM_fft_64_stage_1_0_t343[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t345 = FSM_fft_64_stage_1_0_t329;
    FSM_fft_64_stage_1_0_t345[FSM_fft_64_stage_1_0_t332 * 32 +: 32] = FSM_fft_64_stage_1_0_t344;
    FSM_fft_64_stage_1_0_t346 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001111;
    FSM_fft_64_stage_1_0_t347 = FSM_fft_64_stage_1_0_t346[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t348 = FSM_fft_64_stage_1_0_t347 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t349 = FSM_fft_64_stage_1_0_t348[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t350 = FSM_fft_64_stage_1_0_t349[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t351 = FSM_fft_64_stage_1_0_t345;
    FSM_fft_64_stage_1_0_t351[FSM_fft_64_stage_1_0_t350 * 32 +: 32] = FSM_fft_64_stage_1_0_t336 - FSM_fft_64_stage_1_0_t342;
    FSM_fft_64_stage_1_0_t352 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010000;
    FSM_fft_64_stage_1_0_t353 = FSM_fft_64_stage_1_0_t352[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t354 = FSM_fft_64_stage_1_0_t353[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t355 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010000;
    FSM_fft_64_stage_1_0_t356 = FSM_fft_64_stage_1_0_t355[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t357 = FSM_fft_64_stage_1_0_t356[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t358 = i_data_in_real[FSM_fft_64_stage_1_0_t357 * 32 +: 32];
    FSM_fft_64_stage_1_0_t359 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010000;
    FSM_fft_64_stage_1_0_t360 = FSM_fft_64_stage_1_0_t359[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t361 = FSM_fft_64_stage_1_0_t360 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t362 = FSM_fft_64_stage_1_0_t361[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t363 = FSM_fft_64_stage_1_0_t362[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t364 = i_data_in_real[FSM_fft_64_stage_1_0_t363 * 32 +: 32];
    FSM_fft_64_stage_1_0_t365 = FSM_fft_64_stage_1_0_t358 + FSM_fft_64_stage_1_0_t364;
    FSM_fft_64_stage_1_0_t366 = FSM_fft_64_stage_1_0_t365[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t367 = FSM_fft_64_stage_1_0_t351;
    FSM_fft_64_stage_1_0_t367[FSM_fft_64_stage_1_0_t354 * 32 +: 32] = FSM_fft_64_stage_1_0_t366;
    FSM_fft_64_stage_1_0_t368 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010000;
    FSM_fft_64_stage_1_0_t369 = FSM_fft_64_stage_1_0_t368[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t370 = FSM_fft_64_stage_1_0_t369 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t371 = FSM_fft_64_stage_1_0_t370[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t372 = FSM_fft_64_stage_1_0_t371[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t373 = FSM_fft_64_stage_1_0_t367;
    FSM_fft_64_stage_1_0_t373[FSM_fft_64_stage_1_0_t372 * 32 +: 32] = FSM_fft_64_stage_1_0_t358 - FSM_fft_64_stage_1_0_t364;
    FSM_fft_64_stage_1_0_t374 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010001;
    FSM_fft_64_stage_1_0_t375 = FSM_fft_64_stage_1_0_t374[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t376 = FSM_fft_64_stage_1_0_t375[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t377 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010001;
    FSM_fft_64_stage_1_0_t378 = FSM_fft_64_stage_1_0_t377[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t379 = FSM_fft_64_stage_1_0_t378[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t380 = i_data_in_real[FSM_fft_64_stage_1_0_t379 * 32 +: 32];
    FSM_fft_64_stage_1_0_t381 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010001;
    FSM_fft_64_stage_1_0_t382 = FSM_fft_64_stage_1_0_t381[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t383 = FSM_fft_64_stage_1_0_t382 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t384 = FSM_fft_64_stage_1_0_t383[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t385 = FSM_fft_64_stage_1_0_t384[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t386 = i_data_in_real[FSM_fft_64_stage_1_0_t385 * 32 +: 32];
    FSM_fft_64_stage_1_0_t387 = FSM_fft_64_stage_1_0_t380 + FSM_fft_64_stage_1_0_t386;
    FSM_fft_64_stage_1_0_t388 = FSM_fft_64_stage_1_0_t387[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t389 = FSM_fft_64_stage_1_0_t373;
    FSM_fft_64_stage_1_0_t389[FSM_fft_64_stage_1_0_t376 * 32 +: 32] = FSM_fft_64_stage_1_0_t388;
    FSM_fft_64_stage_1_0_t390 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010001;
    FSM_fft_64_stage_1_0_t391 = FSM_fft_64_stage_1_0_t390[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t392 = FSM_fft_64_stage_1_0_t391 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t393 = FSM_fft_64_stage_1_0_t392[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t394 = FSM_fft_64_stage_1_0_t393[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t395 = FSM_fft_64_stage_1_0_t389;
    FSM_fft_64_stage_1_0_t395[FSM_fft_64_stage_1_0_t394 * 32 +: 32] = FSM_fft_64_stage_1_0_t380 - FSM_fft_64_stage_1_0_t386;
    FSM_fft_64_stage_1_0_t396 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010010;
    FSM_fft_64_stage_1_0_t397 = FSM_fft_64_stage_1_0_t396[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t398 = FSM_fft_64_stage_1_0_t397[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t399 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010010;
    FSM_fft_64_stage_1_0_t400 = FSM_fft_64_stage_1_0_t399[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t401 = FSM_fft_64_stage_1_0_t400[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t402 = i_data_in_real[FSM_fft_64_stage_1_0_t401 * 32 +: 32];
    FSM_fft_64_stage_1_0_t403 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010010;
    FSM_fft_64_stage_1_0_t404 = FSM_fft_64_stage_1_0_t403[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t405 = FSM_fft_64_stage_1_0_t404 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t406 = FSM_fft_64_stage_1_0_t405[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t407 = FSM_fft_64_stage_1_0_t406[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t408 = i_data_in_real[FSM_fft_64_stage_1_0_t407 * 32 +: 32];
    FSM_fft_64_stage_1_0_t409 = FSM_fft_64_stage_1_0_t402 + FSM_fft_64_stage_1_0_t408;
    FSM_fft_64_stage_1_0_t410 = FSM_fft_64_stage_1_0_t409[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t411 = FSM_fft_64_stage_1_0_t395;
    FSM_fft_64_stage_1_0_t411[FSM_fft_64_stage_1_0_t398 * 32 +: 32] = FSM_fft_64_stage_1_0_t410;
    FSM_fft_64_stage_1_0_t412 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010010;
    FSM_fft_64_stage_1_0_t413 = FSM_fft_64_stage_1_0_t412[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t414 = FSM_fft_64_stage_1_0_t413 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t415 = FSM_fft_64_stage_1_0_t414[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t416 = FSM_fft_64_stage_1_0_t415[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t417 = FSM_fft_64_stage_1_0_t411;
    FSM_fft_64_stage_1_0_t417[FSM_fft_64_stage_1_0_t416 * 32 +: 32] = FSM_fft_64_stage_1_0_t402 - FSM_fft_64_stage_1_0_t408;
    FSM_fft_64_stage_1_0_t418 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010011;
    FSM_fft_64_stage_1_0_t419 = FSM_fft_64_stage_1_0_t418[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t420 = FSM_fft_64_stage_1_0_t419[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t421 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010011;
    FSM_fft_64_stage_1_0_t422 = FSM_fft_64_stage_1_0_t421[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t423 = FSM_fft_64_stage_1_0_t422[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t424 = i_data_in_real[FSM_fft_64_stage_1_0_t423 * 32 +: 32];
    FSM_fft_64_stage_1_0_t425 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010011;
    FSM_fft_64_stage_1_0_t426 = FSM_fft_64_stage_1_0_t425[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t427 = FSM_fft_64_stage_1_0_t426 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t428 = FSM_fft_64_stage_1_0_t427[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t429 = FSM_fft_64_stage_1_0_t428[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t430 = i_data_in_real[FSM_fft_64_stage_1_0_t429 * 32 +: 32];
    FSM_fft_64_stage_1_0_t431 = FSM_fft_64_stage_1_0_t424 + FSM_fft_64_stage_1_0_t430;
    FSM_fft_64_stage_1_0_t432 = FSM_fft_64_stage_1_0_t431[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t433 = FSM_fft_64_stage_1_0_t417;
    FSM_fft_64_stage_1_0_t433[FSM_fft_64_stage_1_0_t420 * 32 +: 32] = FSM_fft_64_stage_1_0_t432;
    FSM_fft_64_stage_1_0_t434 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010011;
    FSM_fft_64_stage_1_0_t435 = FSM_fft_64_stage_1_0_t434[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t436 = FSM_fft_64_stage_1_0_t435 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t437 = FSM_fft_64_stage_1_0_t436[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t438 = FSM_fft_64_stage_1_0_t437[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t439 = FSM_fft_64_stage_1_0_t433;
    FSM_fft_64_stage_1_0_t439[FSM_fft_64_stage_1_0_t438 * 32 +: 32] = FSM_fft_64_stage_1_0_t424 - FSM_fft_64_stage_1_0_t430;
    FSM_fft_64_stage_1_0_t440 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010100;
    FSM_fft_64_stage_1_0_t441 = FSM_fft_64_stage_1_0_t440[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t442 = FSM_fft_64_stage_1_0_t441[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t443 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010100;
    FSM_fft_64_stage_1_0_t444 = FSM_fft_64_stage_1_0_t443[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t445 = FSM_fft_64_stage_1_0_t444[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t446 = i_data_in_real[FSM_fft_64_stage_1_0_t445 * 32 +: 32];
    FSM_fft_64_stage_1_0_t447 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010100;
    FSM_fft_64_stage_1_0_t448 = FSM_fft_64_stage_1_0_t447[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t449 = FSM_fft_64_stage_1_0_t448 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t450 = FSM_fft_64_stage_1_0_t449[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t451 = FSM_fft_64_stage_1_0_t450[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t452 = i_data_in_real[FSM_fft_64_stage_1_0_t451 * 32 +: 32];
    FSM_fft_64_stage_1_0_t453 = FSM_fft_64_stage_1_0_t446 + FSM_fft_64_stage_1_0_t452;
    FSM_fft_64_stage_1_0_t454 = FSM_fft_64_stage_1_0_t453[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t455 = FSM_fft_64_stage_1_0_t439;
    FSM_fft_64_stage_1_0_t455[FSM_fft_64_stage_1_0_t442 * 32 +: 32] = FSM_fft_64_stage_1_0_t454;
    FSM_fft_64_stage_1_0_t456 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010100;
    FSM_fft_64_stage_1_0_t457 = FSM_fft_64_stage_1_0_t456[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t458 = FSM_fft_64_stage_1_0_t457 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t459 = FSM_fft_64_stage_1_0_t458[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t460 = FSM_fft_64_stage_1_0_t459[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t461 = FSM_fft_64_stage_1_0_t455;
    FSM_fft_64_stage_1_0_t461[FSM_fft_64_stage_1_0_t460 * 32 +: 32] = FSM_fft_64_stage_1_0_t446 - FSM_fft_64_stage_1_0_t452;
    FSM_fft_64_stage_1_0_t462 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010101;
    FSM_fft_64_stage_1_0_t463 = FSM_fft_64_stage_1_0_t462[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t464 = FSM_fft_64_stage_1_0_t463[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t465 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010101;
    FSM_fft_64_stage_1_0_t466 = FSM_fft_64_stage_1_0_t465[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t467 = FSM_fft_64_stage_1_0_t466[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t468 = i_data_in_real[FSM_fft_64_stage_1_0_t467 * 32 +: 32];
    FSM_fft_64_stage_1_0_t469 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010101;
    FSM_fft_64_stage_1_0_t470 = FSM_fft_64_stage_1_0_t469[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t471 = FSM_fft_64_stage_1_0_t470 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t472 = FSM_fft_64_stage_1_0_t471[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t473 = FSM_fft_64_stage_1_0_t472[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t474 = i_data_in_real[FSM_fft_64_stage_1_0_t473 * 32 +: 32];
    FSM_fft_64_stage_1_0_t475 = FSM_fft_64_stage_1_0_t468 + FSM_fft_64_stage_1_0_t474;
    FSM_fft_64_stage_1_0_t476 = FSM_fft_64_stage_1_0_t475[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t477 = FSM_fft_64_stage_1_0_t461;
    FSM_fft_64_stage_1_0_t477[FSM_fft_64_stage_1_0_t464 * 32 +: 32] = FSM_fft_64_stage_1_0_t476;
    FSM_fft_64_stage_1_0_t478 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010101;
    FSM_fft_64_stage_1_0_t479 = FSM_fft_64_stage_1_0_t478[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t480 = FSM_fft_64_stage_1_0_t479 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t481 = FSM_fft_64_stage_1_0_t480[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t482 = FSM_fft_64_stage_1_0_t481[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t483 = FSM_fft_64_stage_1_0_t477;
    FSM_fft_64_stage_1_0_t483[FSM_fft_64_stage_1_0_t482 * 32 +: 32] = FSM_fft_64_stage_1_0_t468 - FSM_fft_64_stage_1_0_t474;
    FSM_fft_64_stage_1_0_t484 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010110;
    FSM_fft_64_stage_1_0_t485 = FSM_fft_64_stage_1_0_t484[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t486 = FSM_fft_64_stage_1_0_t485[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t487 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010110;
    FSM_fft_64_stage_1_0_t488 = FSM_fft_64_stage_1_0_t487[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t489 = FSM_fft_64_stage_1_0_t488[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t490 = i_data_in_real[FSM_fft_64_stage_1_0_t489 * 32 +: 32];
    FSM_fft_64_stage_1_0_t491 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010110;
    FSM_fft_64_stage_1_0_t492 = FSM_fft_64_stage_1_0_t491[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t493 = FSM_fft_64_stage_1_0_t492 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t494 = FSM_fft_64_stage_1_0_t493[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t495 = FSM_fft_64_stage_1_0_t494[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t496 = i_data_in_real[FSM_fft_64_stage_1_0_t495 * 32 +: 32];
    FSM_fft_64_stage_1_0_t497 = FSM_fft_64_stage_1_0_t490 + FSM_fft_64_stage_1_0_t496;
    FSM_fft_64_stage_1_0_t498 = FSM_fft_64_stage_1_0_t497[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t499 = FSM_fft_64_stage_1_0_t483;
    FSM_fft_64_stage_1_0_t499[FSM_fft_64_stage_1_0_t486 * 32 +: 32] = FSM_fft_64_stage_1_0_t498;
    FSM_fft_64_stage_1_0_t500 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010110;
    FSM_fft_64_stage_1_0_t501 = FSM_fft_64_stage_1_0_t500[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t502 = FSM_fft_64_stage_1_0_t501 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t503 = FSM_fft_64_stage_1_0_t502[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t504 = FSM_fft_64_stage_1_0_t503[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t505 = FSM_fft_64_stage_1_0_t499;
    FSM_fft_64_stage_1_0_t505[FSM_fft_64_stage_1_0_t504 * 32 +: 32] = FSM_fft_64_stage_1_0_t490 - FSM_fft_64_stage_1_0_t496;
    FSM_fft_64_stage_1_0_t506 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010111;
    FSM_fft_64_stage_1_0_t507 = FSM_fft_64_stage_1_0_t506[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t508 = FSM_fft_64_stage_1_0_t507[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t509 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010111;
    FSM_fft_64_stage_1_0_t510 = FSM_fft_64_stage_1_0_t509[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t511 = FSM_fft_64_stage_1_0_t510[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t512 = i_data_in_real[FSM_fft_64_stage_1_0_t511 * 32 +: 32];
    FSM_fft_64_stage_1_0_t513 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010111;
    FSM_fft_64_stage_1_0_t514 = FSM_fft_64_stage_1_0_t513[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t515 = FSM_fft_64_stage_1_0_t514 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t516 = FSM_fft_64_stage_1_0_t515[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t517 = FSM_fft_64_stage_1_0_t516[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t518 = i_data_in_real[FSM_fft_64_stage_1_0_t517 * 32 +: 32];
    FSM_fft_64_stage_1_0_t519 = FSM_fft_64_stage_1_0_t512 + FSM_fft_64_stage_1_0_t518;
    FSM_fft_64_stage_1_0_t520 = FSM_fft_64_stage_1_0_t519[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t521 = FSM_fft_64_stage_1_0_t505;
    FSM_fft_64_stage_1_0_t521[FSM_fft_64_stage_1_0_t508 * 32 +: 32] = FSM_fft_64_stage_1_0_t520;
    FSM_fft_64_stage_1_0_t522 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010111;
    FSM_fft_64_stage_1_0_t523 = FSM_fft_64_stage_1_0_t522[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t524 = FSM_fft_64_stage_1_0_t523 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t525 = FSM_fft_64_stage_1_0_t524[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t526 = FSM_fft_64_stage_1_0_t525[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t527 = FSM_fft_64_stage_1_0_t521;
    FSM_fft_64_stage_1_0_t527[FSM_fft_64_stage_1_0_t526 * 32 +: 32] = FSM_fft_64_stage_1_0_t512 - FSM_fft_64_stage_1_0_t518;
    FSM_fft_64_stage_1_0_t528 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011000;
    FSM_fft_64_stage_1_0_t529 = FSM_fft_64_stage_1_0_t528[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t530 = FSM_fft_64_stage_1_0_t529[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t531 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011000;
    FSM_fft_64_stage_1_0_t532 = FSM_fft_64_stage_1_0_t531[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t533 = FSM_fft_64_stage_1_0_t532[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t534 = i_data_in_real[FSM_fft_64_stage_1_0_t533 * 32 +: 32];
    FSM_fft_64_stage_1_0_t535 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011000;
    FSM_fft_64_stage_1_0_t536 = FSM_fft_64_stage_1_0_t535[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t537 = FSM_fft_64_stage_1_0_t536 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t538 = FSM_fft_64_stage_1_0_t537[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t539 = FSM_fft_64_stage_1_0_t538[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t540 = i_data_in_real[FSM_fft_64_stage_1_0_t539 * 32 +: 32];
    FSM_fft_64_stage_1_0_t541 = FSM_fft_64_stage_1_0_t534 + FSM_fft_64_stage_1_0_t540;
    FSM_fft_64_stage_1_0_t542 = FSM_fft_64_stage_1_0_t541[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t543 = FSM_fft_64_stage_1_0_t527;
    FSM_fft_64_stage_1_0_t543[FSM_fft_64_stage_1_0_t530 * 32 +: 32] = FSM_fft_64_stage_1_0_t542;
    FSM_fft_64_stage_1_0_t544 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011000;
    FSM_fft_64_stage_1_0_t545 = FSM_fft_64_stage_1_0_t544[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t546 = FSM_fft_64_stage_1_0_t545 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t547 = FSM_fft_64_stage_1_0_t546[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t548 = FSM_fft_64_stage_1_0_t547[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t549 = FSM_fft_64_stage_1_0_t543;
    FSM_fft_64_stage_1_0_t549[FSM_fft_64_stage_1_0_t548 * 32 +: 32] = FSM_fft_64_stage_1_0_t534 - FSM_fft_64_stage_1_0_t540;
    FSM_fft_64_stage_1_0_t550 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011001;
    FSM_fft_64_stage_1_0_t551 = FSM_fft_64_stage_1_0_t550[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t552 = FSM_fft_64_stage_1_0_t551[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t553 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011001;
    FSM_fft_64_stage_1_0_t554 = FSM_fft_64_stage_1_0_t553[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t555 = FSM_fft_64_stage_1_0_t554[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t556 = i_data_in_real[FSM_fft_64_stage_1_0_t555 * 32 +: 32];
    FSM_fft_64_stage_1_0_t557 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011001;
    FSM_fft_64_stage_1_0_t558 = FSM_fft_64_stage_1_0_t557[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t559 = FSM_fft_64_stage_1_0_t558 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t560 = FSM_fft_64_stage_1_0_t559[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t561 = FSM_fft_64_stage_1_0_t560[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t562 = i_data_in_real[FSM_fft_64_stage_1_0_t561 * 32 +: 32];
    FSM_fft_64_stage_1_0_t563 = FSM_fft_64_stage_1_0_t556 + FSM_fft_64_stage_1_0_t562;
    FSM_fft_64_stage_1_0_t564 = FSM_fft_64_stage_1_0_t563[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t565 = FSM_fft_64_stage_1_0_t549;
    FSM_fft_64_stage_1_0_t565[FSM_fft_64_stage_1_0_t552 * 32 +: 32] = FSM_fft_64_stage_1_0_t564;
    FSM_fft_64_stage_1_0_t566 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011001;
    FSM_fft_64_stage_1_0_t567 = FSM_fft_64_stage_1_0_t566[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t568 = FSM_fft_64_stage_1_0_t567 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t569 = FSM_fft_64_stage_1_0_t568[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t570 = FSM_fft_64_stage_1_0_t569[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t571 = FSM_fft_64_stage_1_0_t565;
    FSM_fft_64_stage_1_0_t571[FSM_fft_64_stage_1_0_t570 * 32 +: 32] = FSM_fft_64_stage_1_0_t556 - FSM_fft_64_stage_1_0_t562;
    FSM_fft_64_stage_1_0_t572 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011010;
    FSM_fft_64_stage_1_0_t573 = FSM_fft_64_stage_1_0_t572[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t574 = FSM_fft_64_stage_1_0_t573[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t575 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011010;
    FSM_fft_64_stage_1_0_t576 = FSM_fft_64_stage_1_0_t575[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t577 = FSM_fft_64_stage_1_0_t576[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t578 = i_data_in_real[FSM_fft_64_stage_1_0_t577 * 32 +: 32];
    FSM_fft_64_stage_1_0_t579 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011010;
    FSM_fft_64_stage_1_0_t580 = FSM_fft_64_stage_1_0_t579[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t581 = FSM_fft_64_stage_1_0_t580 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t582 = FSM_fft_64_stage_1_0_t581[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t583 = FSM_fft_64_stage_1_0_t582[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t584 = i_data_in_real[FSM_fft_64_stage_1_0_t583 * 32 +: 32];
    FSM_fft_64_stage_1_0_t585 = FSM_fft_64_stage_1_0_t578 + FSM_fft_64_stage_1_0_t584;
    FSM_fft_64_stage_1_0_t586 = FSM_fft_64_stage_1_0_t585[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t587 = FSM_fft_64_stage_1_0_t571;
    FSM_fft_64_stage_1_0_t587[FSM_fft_64_stage_1_0_t574 * 32 +: 32] = FSM_fft_64_stage_1_0_t586;
    FSM_fft_64_stage_1_0_t588 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011010;
    FSM_fft_64_stage_1_0_t589 = FSM_fft_64_stage_1_0_t588[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t590 = FSM_fft_64_stage_1_0_t589 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t591 = FSM_fft_64_stage_1_0_t590[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t592 = FSM_fft_64_stage_1_0_t591[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t593 = FSM_fft_64_stage_1_0_t587;
    FSM_fft_64_stage_1_0_t593[FSM_fft_64_stage_1_0_t592 * 32 +: 32] = FSM_fft_64_stage_1_0_t578 - FSM_fft_64_stage_1_0_t584;
    FSM_fft_64_stage_1_0_t594 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011011;
    FSM_fft_64_stage_1_0_t595 = FSM_fft_64_stage_1_0_t594[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t596 = FSM_fft_64_stage_1_0_t595[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t597 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011011;
    FSM_fft_64_stage_1_0_t598 = FSM_fft_64_stage_1_0_t597[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t599 = FSM_fft_64_stage_1_0_t598[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t600 = i_data_in_real[FSM_fft_64_stage_1_0_t599 * 32 +: 32];
    FSM_fft_64_stage_1_0_t601 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011011;
    FSM_fft_64_stage_1_0_t602 = FSM_fft_64_stage_1_0_t601[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t603 = FSM_fft_64_stage_1_0_t602 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t604 = FSM_fft_64_stage_1_0_t603[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t605 = FSM_fft_64_stage_1_0_t604[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t606 = i_data_in_real[FSM_fft_64_stage_1_0_t605 * 32 +: 32];
    FSM_fft_64_stage_1_0_t607 = FSM_fft_64_stage_1_0_t600 + FSM_fft_64_stage_1_0_t606;
    FSM_fft_64_stage_1_0_t608 = FSM_fft_64_stage_1_0_t607[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t609 = FSM_fft_64_stage_1_0_t593;
    FSM_fft_64_stage_1_0_t609[FSM_fft_64_stage_1_0_t596 * 32 +: 32] = FSM_fft_64_stage_1_0_t608;
    FSM_fft_64_stage_1_0_t610 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011011;
    FSM_fft_64_stage_1_0_t611 = FSM_fft_64_stage_1_0_t610[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t612 = FSM_fft_64_stage_1_0_t611 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t613 = FSM_fft_64_stage_1_0_t612[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t614 = FSM_fft_64_stage_1_0_t613[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t615 = FSM_fft_64_stage_1_0_t609;
    FSM_fft_64_stage_1_0_t615[FSM_fft_64_stage_1_0_t614 * 32 +: 32] = FSM_fft_64_stage_1_0_t600 - FSM_fft_64_stage_1_0_t606;
    FSM_fft_64_stage_1_0_t616 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011100;
    FSM_fft_64_stage_1_0_t617 = FSM_fft_64_stage_1_0_t616[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t618 = FSM_fft_64_stage_1_0_t617[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t619 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011100;
    FSM_fft_64_stage_1_0_t620 = FSM_fft_64_stage_1_0_t619[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t621 = FSM_fft_64_stage_1_0_t620[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t622 = i_data_in_real[FSM_fft_64_stage_1_0_t621 * 32 +: 32];
    FSM_fft_64_stage_1_0_t623 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011100;
    FSM_fft_64_stage_1_0_t624 = FSM_fft_64_stage_1_0_t623[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t625 = FSM_fft_64_stage_1_0_t624 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t626 = FSM_fft_64_stage_1_0_t625[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t627 = FSM_fft_64_stage_1_0_t626[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t628 = i_data_in_real[FSM_fft_64_stage_1_0_t627 * 32 +: 32];
    FSM_fft_64_stage_1_0_t629 = FSM_fft_64_stage_1_0_t622 + FSM_fft_64_stage_1_0_t628;
    FSM_fft_64_stage_1_0_t630 = FSM_fft_64_stage_1_0_t629[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t631 = FSM_fft_64_stage_1_0_t615;
    FSM_fft_64_stage_1_0_t631[FSM_fft_64_stage_1_0_t618 * 32 +: 32] = FSM_fft_64_stage_1_0_t630;
    FSM_fft_64_stage_1_0_t632 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011100;
    FSM_fft_64_stage_1_0_t633 = FSM_fft_64_stage_1_0_t632[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t634 = FSM_fft_64_stage_1_0_t633 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t635 = FSM_fft_64_stage_1_0_t634[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t636 = FSM_fft_64_stage_1_0_t635[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t637 = FSM_fft_64_stage_1_0_t631;
    FSM_fft_64_stage_1_0_t637[FSM_fft_64_stage_1_0_t636 * 32 +: 32] = FSM_fft_64_stage_1_0_t622 - FSM_fft_64_stage_1_0_t628;
    FSM_fft_64_stage_1_0_t638 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011101;
    FSM_fft_64_stage_1_0_t639 = FSM_fft_64_stage_1_0_t638[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t640 = FSM_fft_64_stage_1_0_t639[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t641 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011101;
    FSM_fft_64_stage_1_0_t642 = FSM_fft_64_stage_1_0_t641[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t643 = FSM_fft_64_stage_1_0_t642[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t644 = i_data_in_real[FSM_fft_64_stage_1_0_t643 * 32 +: 32];
    FSM_fft_64_stage_1_0_t645 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011101;
    FSM_fft_64_stage_1_0_t646 = FSM_fft_64_stage_1_0_t645[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t647 = FSM_fft_64_stage_1_0_t646 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t648 = FSM_fft_64_stage_1_0_t647[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t649 = FSM_fft_64_stage_1_0_t648[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t650 = i_data_in_real[FSM_fft_64_stage_1_0_t649 * 32 +: 32];
    FSM_fft_64_stage_1_0_t651 = FSM_fft_64_stage_1_0_t644 + FSM_fft_64_stage_1_0_t650;
    FSM_fft_64_stage_1_0_t652 = FSM_fft_64_stage_1_0_t651[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t653 = FSM_fft_64_stage_1_0_t637;
    FSM_fft_64_stage_1_0_t653[FSM_fft_64_stage_1_0_t640 * 32 +: 32] = FSM_fft_64_stage_1_0_t652;
    FSM_fft_64_stage_1_0_t654 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011101;
    FSM_fft_64_stage_1_0_t655 = FSM_fft_64_stage_1_0_t654[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t656 = FSM_fft_64_stage_1_0_t655 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t657 = FSM_fft_64_stage_1_0_t656[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t658 = FSM_fft_64_stage_1_0_t657[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t659 = FSM_fft_64_stage_1_0_t653;
    FSM_fft_64_stage_1_0_t659[FSM_fft_64_stage_1_0_t658 * 32 +: 32] = FSM_fft_64_stage_1_0_t644 - FSM_fft_64_stage_1_0_t650;
    FSM_fft_64_stage_1_0_t660 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011110;
    FSM_fft_64_stage_1_0_t661 = FSM_fft_64_stage_1_0_t660[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t662 = FSM_fft_64_stage_1_0_t661[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t663 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011110;
    FSM_fft_64_stage_1_0_t664 = FSM_fft_64_stage_1_0_t663[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t665 = FSM_fft_64_stage_1_0_t664[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t666 = i_data_in_real[FSM_fft_64_stage_1_0_t665 * 32 +: 32];
    FSM_fft_64_stage_1_0_t667 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011110;
    FSM_fft_64_stage_1_0_t668 = FSM_fft_64_stage_1_0_t667[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t669 = FSM_fft_64_stage_1_0_t668 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t670 = FSM_fft_64_stage_1_0_t669[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t671 = FSM_fft_64_stage_1_0_t670[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t672 = i_data_in_real[FSM_fft_64_stage_1_0_t671 * 32 +: 32];
    FSM_fft_64_stage_1_0_t673 = FSM_fft_64_stage_1_0_t666 + FSM_fft_64_stage_1_0_t672;
    FSM_fft_64_stage_1_0_t674 = FSM_fft_64_stage_1_0_t673[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t675 = FSM_fft_64_stage_1_0_t659;
    FSM_fft_64_stage_1_0_t675[FSM_fft_64_stage_1_0_t662 * 32 +: 32] = FSM_fft_64_stage_1_0_t674;
    FSM_fft_64_stage_1_0_t676 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011110;
    FSM_fft_64_stage_1_0_t677 = FSM_fft_64_stage_1_0_t676[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t678 = FSM_fft_64_stage_1_0_t677 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t679 = FSM_fft_64_stage_1_0_t678[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t680 = FSM_fft_64_stage_1_0_t679[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t681 = FSM_fft_64_stage_1_0_t675;
    FSM_fft_64_stage_1_0_t681[FSM_fft_64_stage_1_0_t680 * 32 +: 32] = FSM_fft_64_stage_1_0_t666 - FSM_fft_64_stage_1_0_t672;
    FSM_fft_64_stage_1_0_t682 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011111;
    FSM_fft_64_stage_1_0_t683 = FSM_fft_64_stage_1_0_t682[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t684 = FSM_fft_64_stage_1_0_t683[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t685 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011111;
    FSM_fft_64_stage_1_0_t686 = FSM_fft_64_stage_1_0_t685[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t687 = FSM_fft_64_stage_1_0_t686[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t688 = i_data_in_real[FSM_fft_64_stage_1_0_t687 * 32 +: 32];
    FSM_fft_64_stage_1_0_t689 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011111;
    FSM_fft_64_stage_1_0_t690 = FSM_fft_64_stage_1_0_t689[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t691 = FSM_fft_64_stage_1_0_t690 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t692 = FSM_fft_64_stage_1_0_t691[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t693 = FSM_fft_64_stage_1_0_t692[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t694 = i_data_in_real[FSM_fft_64_stage_1_0_t693 * 32 +: 32];
    FSM_fft_64_stage_1_0_t695 = FSM_fft_64_stage_1_0_t688 + FSM_fft_64_stage_1_0_t694;
    FSM_fft_64_stage_1_0_t696 = FSM_fft_64_stage_1_0_t695[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t697 = FSM_fft_64_stage_1_0_t681;
    FSM_fft_64_stage_1_0_t697[FSM_fft_64_stage_1_0_t684 * 32 +: 32] = FSM_fft_64_stage_1_0_t696;
    FSM_fft_64_stage_1_0_t698 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011111;
    FSM_fft_64_stage_1_0_t699 = FSM_fft_64_stage_1_0_t698[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t700 = FSM_fft_64_stage_1_0_t699 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t701 = FSM_fft_64_stage_1_0_t700[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t702 = FSM_fft_64_stage_1_0_t701[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t703 = FSM_fft_64_stage_1_0_t697;
    FSM_fft_64_stage_1_0_t703[FSM_fft_64_stage_1_0_t702 * 32 +: 32] = FSM_fft_64_stage_1_0_t688 - FSM_fft_64_stage_1_0_t694;
    FSM_fft_64_stage_1_0_t704 = 32'b00000000000000000000000000000010 * 32'b0;
    FSM_fft_64_stage_1_0_t705 = FSM_fft_64_stage_1_0_t704[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t706 = FSM_fft_64_stage_1_0_t705[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t707 = 32'b00000000000000000000000000000010 * 32'b0;
    FSM_fft_64_stage_1_0_t708 = FSM_fft_64_stage_1_0_t707[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t709 = FSM_fft_64_stage_1_0_t708[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t710 = i_data_in_imag[FSM_fft_64_stage_1_0_t709 * 32 +: 32];
    FSM_fft_64_stage_1_0_t711 = 32'b00000000000000000000000000000010 * 32'b0;
    FSM_fft_64_stage_1_0_t712 = FSM_fft_64_stage_1_0_t711[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t713 = FSM_fft_64_stage_1_0_t712 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t714 = FSM_fft_64_stage_1_0_t713[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t715 = FSM_fft_64_stage_1_0_t714[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t716 = i_data_in_imag[FSM_fft_64_stage_1_0_t715 * 32 +: 32];
    FSM_fft_64_stage_1_0_t717 = FSM_fft_64_stage_1_0_t710 + FSM_fft_64_stage_1_0_t716;
    FSM_fft_64_stage_1_0_t718 = FSM_fft_64_stage_1_0_t717[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t719 = 2048'b0;
    FSM_fft_64_stage_1_0_t719[FSM_fft_64_stage_1_0_t706 * 32 +: 32] = FSM_fft_64_stage_1_0_t718;
    FSM_fft_64_stage_1_0_t720 = 32'b00000000000000000000000000000010 * 32'b0;
    FSM_fft_64_stage_1_0_t721 = FSM_fft_64_stage_1_0_t720[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t722 = FSM_fft_64_stage_1_0_t721 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t723 = FSM_fft_64_stage_1_0_t722[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t724 = FSM_fft_64_stage_1_0_t723[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t725 = FSM_fft_64_stage_1_0_t719;
    FSM_fft_64_stage_1_0_t725[FSM_fft_64_stage_1_0_t724 * 32 +: 32] = FSM_fft_64_stage_1_0_t710 - FSM_fft_64_stage_1_0_t716;
    FSM_fft_64_stage_1_0_t726 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t727 = FSM_fft_64_stage_1_0_t726[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t728 = FSM_fft_64_stage_1_0_t727[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t729 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t730 = FSM_fft_64_stage_1_0_t729[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t731 = FSM_fft_64_stage_1_0_t730[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t732 = i_data_in_imag[FSM_fft_64_stage_1_0_t731 * 32 +: 32];
    FSM_fft_64_stage_1_0_t733 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t734 = FSM_fft_64_stage_1_0_t733[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t735 = FSM_fft_64_stage_1_0_t734 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t736 = FSM_fft_64_stage_1_0_t735[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t737 = FSM_fft_64_stage_1_0_t736[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t738 = i_data_in_imag[FSM_fft_64_stage_1_0_t737 * 32 +: 32];
    FSM_fft_64_stage_1_0_t739 = FSM_fft_64_stage_1_0_t732 + FSM_fft_64_stage_1_0_t738;
    FSM_fft_64_stage_1_0_t740 = FSM_fft_64_stage_1_0_t739[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t741 = FSM_fft_64_stage_1_0_t725;
    FSM_fft_64_stage_1_0_t741[FSM_fft_64_stage_1_0_t728 * 32 +: 32] = FSM_fft_64_stage_1_0_t740;
    FSM_fft_64_stage_1_0_t742 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t743 = FSM_fft_64_stage_1_0_t742[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t744 = FSM_fft_64_stage_1_0_t743 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t745 = FSM_fft_64_stage_1_0_t744[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t746 = FSM_fft_64_stage_1_0_t745[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t747 = FSM_fft_64_stage_1_0_t741;
    FSM_fft_64_stage_1_0_t747[FSM_fft_64_stage_1_0_t746 * 32 +: 32] = FSM_fft_64_stage_1_0_t732 - FSM_fft_64_stage_1_0_t738;
    FSM_fft_64_stage_1_0_t748 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_1_0_t749 = FSM_fft_64_stage_1_0_t748[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t750 = FSM_fft_64_stage_1_0_t749[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t751 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_1_0_t752 = FSM_fft_64_stage_1_0_t751[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t753 = FSM_fft_64_stage_1_0_t752[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t754 = i_data_in_imag[FSM_fft_64_stage_1_0_t753 * 32 +: 32];
    FSM_fft_64_stage_1_0_t755 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_1_0_t756 = FSM_fft_64_stage_1_0_t755[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t757 = FSM_fft_64_stage_1_0_t756 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t758 = FSM_fft_64_stage_1_0_t757[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t759 = FSM_fft_64_stage_1_0_t758[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t760 = i_data_in_imag[FSM_fft_64_stage_1_0_t759 * 32 +: 32];
    FSM_fft_64_stage_1_0_t761 = FSM_fft_64_stage_1_0_t754 + FSM_fft_64_stage_1_0_t760;
    FSM_fft_64_stage_1_0_t762 = FSM_fft_64_stage_1_0_t761[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t763 = FSM_fft_64_stage_1_0_t747;
    FSM_fft_64_stage_1_0_t763[FSM_fft_64_stage_1_0_t750 * 32 +: 32] = FSM_fft_64_stage_1_0_t762;
    FSM_fft_64_stage_1_0_t764 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_1_0_t765 = FSM_fft_64_stage_1_0_t764[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t766 = FSM_fft_64_stage_1_0_t765 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t767 = FSM_fft_64_stage_1_0_t766[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t768 = FSM_fft_64_stage_1_0_t767[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t769 = FSM_fft_64_stage_1_0_t763;
    FSM_fft_64_stage_1_0_t769[FSM_fft_64_stage_1_0_t768 * 32 +: 32] = FSM_fft_64_stage_1_0_t754 - FSM_fft_64_stage_1_0_t760;
    FSM_fft_64_stage_1_0_t770 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_1_0_t771 = FSM_fft_64_stage_1_0_t770[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t772 = FSM_fft_64_stage_1_0_t771[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t773 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_1_0_t774 = FSM_fft_64_stage_1_0_t773[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t775 = FSM_fft_64_stage_1_0_t774[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t776 = i_data_in_imag[FSM_fft_64_stage_1_0_t775 * 32 +: 32];
    FSM_fft_64_stage_1_0_t777 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_1_0_t778 = FSM_fft_64_stage_1_0_t777[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t779 = FSM_fft_64_stage_1_0_t778 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t780 = FSM_fft_64_stage_1_0_t779[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t781 = FSM_fft_64_stage_1_0_t780[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t782 = i_data_in_imag[FSM_fft_64_stage_1_0_t781 * 32 +: 32];
    FSM_fft_64_stage_1_0_t783 = FSM_fft_64_stage_1_0_t776 + FSM_fft_64_stage_1_0_t782;
    FSM_fft_64_stage_1_0_t784 = FSM_fft_64_stage_1_0_t783[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t785 = FSM_fft_64_stage_1_0_t769;
    FSM_fft_64_stage_1_0_t785[FSM_fft_64_stage_1_0_t772 * 32 +: 32] = FSM_fft_64_stage_1_0_t784;
    FSM_fft_64_stage_1_0_t786 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_1_0_t787 = FSM_fft_64_stage_1_0_t786[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t788 = FSM_fft_64_stage_1_0_t787 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t789 = FSM_fft_64_stage_1_0_t788[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t790 = FSM_fft_64_stage_1_0_t789[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t791 = FSM_fft_64_stage_1_0_t785;
    FSM_fft_64_stage_1_0_t791[FSM_fft_64_stage_1_0_t790 * 32 +: 32] = FSM_fft_64_stage_1_0_t776 - FSM_fft_64_stage_1_0_t782;
    FSM_fft_64_stage_1_0_t792 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000100;
    FSM_fft_64_stage_1_0_t793 = FSM_fft_64_stage_1_0_t792[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t794 = FSM_fft_64_stage_1_0_t793[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t795 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000100;
    FSM_fft_64_stage_1_0_t796 = FSM_fft_64_stage_1_0_t795[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t797 = FSM_fft_64_stage_1_0_t796[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t798 = i_data_in_imag[FSM_fft_64_stage_1_0_t797 * 32 +: 32];
    FSM_fft_64_stage_1_0_t799 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000100;
    FSM_fft_64_stage_1_0_t800 = FSM_fft_64_stage_1_0_t799[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t801 = FSM_fft_64_stage_1_0_t800 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t802 = FSM_fft_64_stage_1_0_t801[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t803 = FSM_fft_64_stage_1_0_t802[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t804 = i_data_in_imag[FSM_fft_64_stage_1_0_t803 * 32 +: 32];
    FSM_fft_64_stage_1_0_t805 = FSM_fft_64_stage_1_0_t798 + FSM_fft_64_stage_1_0_t804;
    FSM_fft_64_stage_1_0_t806 = FSM_fft_64_stage_1_0_t805[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t807 = FSM_fft_64_stage_1_0_t791;
    FSM_fft_64_stage_1_0_t807[FSM_fft_64_stage_1_0_t794 * 32 +: 32] = FSM_fft_64_stage_1_0_t806;
    FSM_fft_64_stage_1_0_t808 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000100;
    FSM_fft_64_stage_1_0_t809 = FSM_fft_64_stage_1_0_t808[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t810 = FSM_fft_64_stage_1_0_t809 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t811 = FSM_fft_64_stage_1_0_t810[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t812 = FSM_fft_64_stage_1_0_t811[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t813 = FSM_fft_64_stage_1_0_t807;
    FSM_fft_64_stage_1_0_t813[FSM_fft_64_stage_1_0_t812 * 32 +: 32] = FSM_fft_64_stage_1_0_t798 - FSM_fft_64_stage_1_0_t804;
    FSM_fft_64_stage_1_0_t814 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000101;
    FSM_fft_64_stage_1_0_t815 = FSM_fft_64_stage_1_0_t814[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t816 = FSM_fft_64_stage_1_0_t815[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t817 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000101;
    FSM_fft_64_stage_1_0_t818 = FSM_fft_64_stage_1_0_t817[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t819 = FSM_fft_64_stage_1_0_t818[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t820 = i_data_in_imag[FSM_fft_64_stage_1_0_t819 * 32 +: 32];
    FSM_fft_64_stage_1_0_t821 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000101;
    FSM_fft_64_stage_1_0_t822 = FSM_fft_64_stage_1_0_t821[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t823 = FSM_fft_64_stage_1_0_t822 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t824 = FSM_fft_64_stage_1_0_t823[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t825 = FSM_fft_64_stage_1_0_t824[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t826 = i_data_in_imag[FSM_fft_64_stage_1_0_t825 * 32 +: 32];
    FSM_fft_64_stage_1_0_t827 = FSM_fft_64_stage_1_0_t820 + FSM_fft_64_stage_1_0_t826;
    FSM_fft_64_stage_1_0_t828 = FSM_fft_64_stage_1_0_t827[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t829 = FSM_fft_64_stage_1_0_t813;
    FSM_fft_64_stage_1_0_t829[FSM_fft_64_stage_1_0_t816 * 32 +: 32] = FSM_fft_64_stage_1_0_t828;
    FSM_fft_64_stage_1_0_t830 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000101;
    FSM_fft_64_stage_1_0_t831 = FSM_fft_64_stage_1_0_t830[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t832 = FSM_fft_64_stage_1_0_t831 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t833 = FSM_fft_64_stage_1_0_t832[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t834 = FSM_fft_64_stage_1_0_t833[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t835 = FSM_fft_64_stage_1_0_t829;
    FSM_fft_64_stage_1_0_t835[FSM_fft_64_stage_1_0_t834 * 32 +: 32] = FSM_fft_64_stage_1_0_t820 - FSM_fft_64_stage_1_0_t826;
    FSM_fft_64_stage_1_0_t836 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000110;
    FSM_fft_64_stage_1_0_t837 = FSM_fft_64_stage_1_0_t836[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t838 = FSM_fft_64_stage_1_0_t837[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t839 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000110;
    FSM_fft_64_stage_1_0_t840 = FSM_fft_64_stage_1_0_t839[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t841 = FSM_fft_64_stage_1_0_t840[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t842 = i_data_in_imag[FSM_fft_64_stage_1_0_t841 * 32 +: 32];
    FSM_fft_64_stage_1_0_t843 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000110;
    FSM_fft_64_stage_1_0_t844 = FSM_fft_64_stage_1_0_t843[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t845 = FSM_fft_64_stage_1_0_t844 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t846 = FSM_fft_64_stage_1_0_t845[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t847 = FSM_fft_64_stage_1_0_t846[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t848 = i_data_in_imag[FSM_fft_64_stage_1_0_t847 * 32 +: 32];
    FSM_fft_64_stage_1_0_t849 = FSM_fft_64_stage_1_0_t842 + FSM_fft_64_stage_1_0_t848;
    FSM_fft_64_stage_1_0_t850 = FSM_fft_64_stage_1_0_t849[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t851 = FSM_fft_64_stage_1_0_t835;
    FSM_fft_64_stage_1_0_t851[FSM_fft_64_stage_1_0_t838 * 32 +: 32] = FSM_fft_64_stage_1_0_t850;
    FSM_fft_64_stage_1_0_t852 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000110;
    FSM_fft_64_stage_1_0_t853 = FSM_fft_64_stage_1_0_t852[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t854 = FSM_fft_64_stage_1_0_t853 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t855 = FSM_fft_64_stage_1_0_t854[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t856 = FSM_fft_64_stage_1_0_t855[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t857 = FSM_fft_64_stage_1_0_t851;
    FSM_fft_64_stage_1_0_t857[FSM_fft_64_stage_1_0_t856 * 32 +: 32] = FSM_fft_64_stage_1_0_t842 - FSM_fft_64_stage_1_0_t848;
    FSM_fft_64_stage_1_0_t858 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000111;
    FSM_fft_64_stage_1_0_t859 = FSM_fft_64_stage_1_0_t858[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t860 = FSM_fft_64_stage_1_0_t859[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t861 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000111;
    FSM_fft_64_stage_1_0_t862 = FSM_fft_64_stage_1_0_t861[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t863 = FSM_fft_64_stage_1_0_t862[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t864 = i_data_in_imag[FSM_fft_64_stage_1_0_t863 * 32 +: 32];
    FSM_fft_64_stage_1_0_t865 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000111;
    FSM_fft_64_stage_1_0_t866 = FSM_fft_64_stage_1_0_t865[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t867 = FSM_fft_64_stage_1_0_t866 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t868 = FSM_fft_64_stage_1_0_t867[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t869 = FSM_fft_64_stage_1_0_t868[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t870 = i_data_in_imag[FSM_fft_64_stage_1_0_t869 * 32 +: 32];
    FSM_fft_64_stage_1_0_t871 = FSM_fft_64_stage_1_0_t864 + FSM_fft_64_stage_1_0_t870;
    FSM_fft_64_stage_1_0_t872 = FSM_fft_64_stage_1_0_t871[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t873 = FSM_fft_64_stage_1_0_t857;
    FSM_fft_64_stage_1_0_t873[FSM_fft_64_stage_1_0_t860 * 32 +: 32] = FSM_fft_64_stage_1_0_t872;
    FSM_fft_64_stage_1_0_t874 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000111;
    FSM_fft_64_stage_1_0_t875 = FSM_fft_64_stage_1_0_t874[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t876 = FSM_fft_64_stage_1_0_t875 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t877 = FSM_fft_64_stage_1_0_t876[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t878 = FSM_fft_64_stage_1_0_t877[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t879 = FSM_fft_64_stage_1_0_t873;
    FSM_fft_64_stage_1_0_t879[FSM_fft_64_stage_1_0_t878 * 32 +: 32] = FSM_fft_64_stage_1_0_t864 - FSM_fft_64_stage_1_0_t870;
    FSM_fft_64_stage_1_0_t880 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001000;
    FSM_fft_64_stage_1_0_t881 = FSM_fft_64_stage_1_0_t880[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t882 = FSM_fft_64_stage_1_0_t881[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t883 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001000;
    FSM_fft_64_stage_1_0_t884 = FSM_fft_64_stage_1_0_t883[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t885 = FSM_fft_64_stage_1_0_t884[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t886 = i_data_in_imag[FSM_fft_64_stage_1_0_t885 * 32 +: 32];
    FSM_fft_64_stage_1_0_t887 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001000;
    FSM_fft_64_stage_1_0_t888 = FSM_fft_64_stage_1_0_t887[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t889 = FSM_fft_64_stage_1_0_t888 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t890 = FSM_fft_64_stage_1_0_t889[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t891 = FSM_fft_64_stage_1_0_t890[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t892 = i_data_in_imag[FSM_fft_64_stage_1_0_t891 * 32 +: 32];
    FSM_fft_64_stage_1_0_t893 = FSM_fft_64_stage_1_0_t886 + FSM_fft_64_stage_1_0_t892;
    FSM_fft_64_stage_1_0_t894 = FSM_fft_64_stage_1_0_t893[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t895 = FSM_fft_64_stage_1_0_t879;
    FSM_fft_64_stage_1_0_t895[FSM_fft_64_stage_1_0_t882 * 32 +: 32] = FSM_fft_64_stage_1_0_t894;
    FSM_fft_64_stage_1_0_t896 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001000;
    FSM_fft_64_stage_1_0_t897 = FSM_fft_64_stage_1_0_t896[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t898 = FSM_fft_64_stage_1_0_t897 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t899 = FSM_fft_64_stage_1_0_t898[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t900 = FSM_fft_64_stage_1_0_t899[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t901 = FSM_fft_64_stage_1_0_t895;
    FSM_fft_64_stage_1_0_t901[FSM_fft_64_stage_1_0_t900 * 32 +: 32] = FSM_fft_64_stage_1_0_t886 - FSM_fft_64_stage_1_0_t892;
    FSM_fft_64_stage_1_0_t902 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001001;
    FSM_fft_64_stage_1_0_t903 = FSM_fft_64_stage_1_0_t902[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t904 = FSM_fft_64_stage_1_0_t903[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t905 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001001;
    FSM_fft_64_stage_1_0_t906 = FSM_fft_64_stage_1_0_t905[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t907 = FSM_fft_64_stage_1_0_t906[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t908 = i_data_in_imag[FSM_fft_64_stage_1_0_t907 * 32 +: 32];
    FSM_fft_64_stage_1_0_t909 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001001;
    FSM_fft_64_stage_1_0_t910 = FSM_fft_64_stage_1_0_t909[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t911 = FSM_fft_64_stage_1_0_t910 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t912 = FSM_fft_64_stage_1_0_t911[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t913 = FSM_fft_64_stage_1_0_t912[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t914 = i_data_in_imag[FSM_fft_64_stage_1_0_t913 * 32 +: 32];
    FSM_fft_64_stage_1_0_t915 = FSM_fft_64_stage_1_0_t908 + FSM_fft_64_stage_1_0_t914;
    FSM_fft_64_stage_1_0_t916 = FSM_fft_64_stage_1_0_t915[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t917 = FSM_fft_64_stage_1_0_t901;
    FSM_fft_64_stage_1_0_t917[FSM_fft_64_stage_1_0_t904 * 32 +: 32] = FSM_fft_64_stage_1_0_t916;
    FSM_fft_64_stage_1_0_t918 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001001;
    FSM_fft_64_stage_1_0_t919 = FSM_fft_64_stage_1_0_t918[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t920 = FSM_fft_64_stage_1_0_t919 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t921 = FSM_fft_64_stage_1_0_t920[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t922 = FSM_fft_64_stage_1_0_t921[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t923 = FSM_fft_64_stage_1_0_t917;
    FSM_fft_64_stage_1_0_t923[FSM_fft_64_stage_1_0_t922 * 32 +: 32] = FSM_fft_64_stage_1_0_t908 - FSM_fft_64_stage_1_0_t914;
    FSM_fft_64_stage_1_0_t924 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001010;
    FSM_fft_64_stage_1_0_t925 = FSM_fft_64_stage_1_0_t924[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t926 = FSM_fft_64_stage_1_0_t925[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t927 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001010;
    FSM_fft_64_stage_1_0_t928 = FSM_fft_64_stage_1_0_t927[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t929 = FSM_fft_64_stage_1_0_t928[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t930 = i_data_in_imag[FSM_fft_64_stage_1_0_t929 * 32 +: 32];
    FSM_fft_64_stage_1_0_t931 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001010;
    FSM_fft_64_stage_1_0_t932 = FSM_fft_64_stage_1_0_t931[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t933 = FSM_fft_64_stage_1_0_t932 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t934 = FSM_fft_64_stage_1_0_t933[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t935 = FSM_fft_64_stage_1_0_t934[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t936 = i_data_in_imag[FSM_fft_64_stage_1_0_t935 * 32 +: 32];
    FSM_fft_64_stage_1_0_t937 = FSM_fft_64_stage_1_0_t930 + FSM_fft_64_stage_1_0_t936;
    FSM_fft_64_stage_1_0_t938 = FSM_fft_64_stage_1_0_t937[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t939 = FSM_fft_64_stage_1_0_t923;
    FSM_fft_64_stage_1_0_t939[FSM_fft_64_stage_1_0_t926 * 32 +: 32] = FSM_fft_64_stage_1_0_t938;
    FSM_fft_64_stage_1_0_t940 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001010;
    FSM_fft_64_stage_1_0_t941 = FSM_fft_64_stage_1_0_t940[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t942 = FSM_fft_64_stage_1_0_t941 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t943 = FSM_fft_64_stage_1_0_t942[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t944 = FSM_fft_64_stage_1_0_t943[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t945 = FSM_fft_64_stage_1_0_t939;
    FSM_fft_64_stage_1_0_t945[FSM_fft_64_stage_1_0_t944 * 32 +: 32] = FSM_fft_64_stage_1_0_t930 - FSM_fft_64_stage_1_0_t936;
    FSM_fft_64_stage_1_0_t946 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001011;
    FSM_fft_64_stage_1_0_t947 = FSM_fft_64_stage_1_0_t946[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t948 = FSM_fft_64_stage_1_0_t947[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t949 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001011;
    FSM_fft_64_stage_1_0_t950 = FSM_fft_64_stage_1_0_t949[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t951 = FSM_fft_64_stage_1_0_t950[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t952 = i_data_in_imag[FSM_fft_64_stage_1_0_t951 * 32 +: 32];
    FSM_fft_64_stage_1_0_t953 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001011;
    FSM_fft_64_stage_1_0_t954 = FSM_fft_64_stage_1_0_t953[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t955 = FSM_fft_64_stage_1_0_t954 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t956 = FSM_fft_64_stage_1_0_t955[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t957 = FSM_fft_64_stage_1_0_t956[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t958 = i_data_in_imag[FSM_fft_64_stage_1_0_t957 * 32 +: 32];
    FSM_fft_64_stage_1_0_t959 = FSM_fft_64_stage_1_0_t952 + FSM_fft_64_stage_1_0_t958;
    FSM_fft_64_stage_1_0_t960 = FSM_fft_64_stage_1_0_t959[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t961 = FSM_fft_64_stage_1_0_t945;
    FSM_fft_64_stage_1_0_t961[FSM_fft_64_stage_1_0_t948 * 32 +: 32] = FSM_fft_64_stage_1_0_t960;
    FSM_fft_64_stage_1_0_t962 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001011;
    FSM_fft_64_stage_1_0_t963 = FSM_fft_64_stage_1_0_t962[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t964 = FSM_fft_64_stage_1_0_t963 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t965 = FSM_fft_64_stage_1_0_t964[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t966 = FSM_fft_64_stage_1_0_t965[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t967 = FSM_fft_64_stage_1_0_t961;
    FSM_fft_64_stage_1_0_t967[FSM_fft_64_stage_1_0_t966 * 32 +: 32] = FSM_fft_64_stage_1_0_t952 - FSM_fft_64_stage_1_0_t958;
    FSM_fft_64_stage_1_0_t968 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001100;
    FSM_fft_64_stage_1_0_t969 = FSM_fft_64_stage_1_0_t968[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t970 = FSM_fft_64_stage_1_0_t969[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t971 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001100;
    FSM_fft_64_stage_1_0_t972 = FSM_fft_64_stage_1_0_t971[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t973 = FSM_fft_64_stage_1_0_t972[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t974 = i_data_in_imag[FSM_fft_64_stage_1_0_t973 * 32 +: 32];
    FSM_fft_64_stage_1_0_t975 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001100;
    FSM_fft_64_stage_1_0_t976 = FSM_fft_64_stage_1_0_t975[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t977 = FSM_fft_64_stage_1_0_t976 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t978 = FSM_fft_64_stage_1_0_t977[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t979 = FSM_fft_64_stage_1_0_t978[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t980 = i_data_in_imag[FSM_fft_64_stage_1_0_t979 * 32 +: 32];
    FSM_fft_64_stage_1_0_t981 = FSM_fft_64_stage_1_0_t974 + FSM_fft_64_stage_1_0_t980;
    FSM_fft_64_stage_1_0_t982 = FSM_fft_64_stage_1_0_t981[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t983 = FSM_fft_64_stage_1_0_t967;
    FSM_fft_64_stage_1_0_t983[FSM_fft_64_stage_1_0_t970 * 32 +: 32] = FSM_fft_64_stage_1_0_t982;
    FSM_fft_64_stage_1_0_t984 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001100;
    FSM_fft_64_stage_1_0_t985 = FSM_fft_64_stage_1_0_t984[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t986 = FSM_fft_64_stage_1_0_t985 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t987 = FSM_fft_64_stage_1_0_t986[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t988 = FSM_fft_64_stage_1_0_t987[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t989 = FSM_fft_64_stage_1_0_t983;
    FSM_fft_64_stage_1_0_t989[FSM_fft_64_stage_1_0_t988 * 32 +: 32] = FSM_fft_64_stage_1_0_t974 - FSM_fft_64_stage_1_0_t980;
    FSM_fft_64_stage_1_0_t990 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001101;
    FSM_fft_64_stage_1_0_t991 = FSM_fft_64_stage_1_0_t990[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t992 = FSM_fft_64_stage_1_0_t991[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t993 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001101;
    FSM_fft_64_stage_1_0_t994 = FSM_fft_64_stage_1_0_t993[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t995 = FSM_fft_64_stage_1_0_t994[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t996 = i_data_in_imag[FSM_fft_64_stage_1_0_t995 * 32 +: 32];
    FSM_fft_64_stage_1_0_t997 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001101;
    FSM_fft_64_stage_1_0_t998 = FSM_fft_64_stage_1_0_t997[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t999 = FSM_fft_64_stage_1_0_t998 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1000 = FSM_fft_64_stage_1_0_t999[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1001 = FSM_fft_64_stage_1_0_t1000[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1002 = i_data_in_imag[FSM_fft_64_stage_1_0_t1001 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1003 = FSM_fft_64_stage_1_0_t996 + FSM_fft_64_stage_1_0_t1002;
    FSM_fft_64_stage_1_0_t1004 = FSM_fft_64_stage_1_0_t1003[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1005 = FSM_fft_64_stage_1_0_t989;
    FSM_fft_64_stage_1_0_t1005[FSM_fft_64_stage_1_0_t992 * 32 +: 32] = FSM_fft_64_stage_1_0_t1004;
    FSM_fft_64_stage_1_0_t1006 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001101;
    FSM_fft_64_stage_1_0_t1007 = FSM_fft_64_stage_1_0_t1006[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1008 = FSM_fft_64_stage_1_0_t1007 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1009 = FSM_fft_64_stage_1_0_t1008[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1010 = FSM_fft_64_stage_1_0_t1009[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1011 = FSM_fft_64_stage_1_0_t1005;
    FSM_fft_64_stage_1_0_t1011[FSM_fft_64_stage_1_0_t1010 * 32 +: 32] = FSM_fft_64_stage_1_0_t996 - FSM_fft_64_stage_1_0_t1002;
    FSM_fft_64_stage_1_0_t1012 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001110;
    FSM_fft_64_stage_1_0_t1013 = FSM_fft_64_stage_1_0_t1012[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1014 = FSM_fft_64_stage_1_0_t1013[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1015 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001110;
    FSM_fft_64_stage_1_0_t1016 = FSM_fft_64_stage_1_0_t1015[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1017 = FSM_fft_64_stage_1_0_t1016[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1018 = i_data_in_imag[FSM_fft_64_stage_1_0_t1017 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1019 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001110;
    FSM_fft_64_stage_1_0_t1020 = FSM_fft_64_stage_1_0_t1019[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1021 = FSM_fft_64_stage_1_0_t1020 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1022 = FSM_fft_64_stage_1_0_t1021[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1023 = FSM_fft_64_stage_1_0_t1022[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1024 = i_data_in_imag[FSM_fft_64_stage_1_0_t1023 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1025 = FSM_fft_64_stage_1_0_t1018 + FSM_fft_64_stage_1_0_t1024;
    FSM_fft_64_stage_1_0_t1026 = FSM_fft_64_stage_1_0_t1025[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1027 = FSM_fft_64_stage_1_0_t1011;
    FSM_fft_64_stage_1_0_t1027[FSM_fft_64_stage_1_0_t1014 * 32 +: 32] = FSM_fft_64_stage_1_0_t1026;
    FSM_fft_64_stage_1_0_t1028 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001110;
    FSM_fft_64_stage_1_0_t1029 = FSM_fft_64_stage_1_0_t1028[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1030 = FSM_fft_64_stage_1_0_t1029 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1031 = FSM_fft_64_stage_1_0_t1030[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1032 = FSM_fft_64_stage_1_0_t1031[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1033 = FSM_fft_64_stage_1_0_t1027;
    FSM_fft_64_stage_1_0_t1033[FSM_fft_64_stage_1_0_t1032 * 32 +: 32] = FSM_fft_64_stage_1_0_t1018 - FSM_fft_64_stage_1_0_t1024;
    FSM_fft_64_stage_1_0_t1034 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001111;
    FSM_fft_64_stage_1_0_t1035 = FSM_fft_64_stage_1_0_t1034[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1036 = FSM_fft_64_stage_1_0_t1035[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1037 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001111;
    FSM_fft_64_stage_1_0_t1038 = FSM_fft_64_stage_1_0_t1037[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1039 = FSM_fft_64_stage_1_0_t1038[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1040 = i_data_in_imag[FSM_fft_64_stage_1_0_t1039 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1041 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001111;
    FSM_fft_64_stage_1_0_t1042 = FSM_fft_64_stage_1_0_t1041[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1043 = FSM_fft_64_stage_1_0_t1042 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1044 = FSM_fft_64_stage_1_0_t1043[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1045 = FSM_fft_64_stage_1_0_t1044[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1046 = i_data_in_imag[FSM_fft_64_stage_1_0_t1045 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1047 = FSM_fft_64_stage_1_0_t1040 + FSM_fft_64_stage_1_0_t1046;
    FSM_fft_64_stage_1_0_t1048 = FSM_fft_64_stage_1_0_t1047[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1049 = FSM_fft_64_stage_1_0_t1033;
    FSM_fft_64_stage_1_0_t1049[FSM_fft_64_stage_1_0_t1036 * 32 +: 32] = FSM_fft_64_stage_1_0_t1048;
    FSM_fft_64_stage_1_0_t1050 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001111;
    FSM_fft_64_stage_1_0_t1051 = FSM_fft_64_stage_1_0_t1050[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1052 = FSM_fft_64_stage_1_0_t1051 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1053 = FSM_fft_64_stage_1_0_t1052[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1054 = FSM_fft_64_stage_1_0_t1053[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1055 = FSM_fft_64_stage_1_0_t1049;
    FSM_fft_64_stage_1_0_t1055[FSM_fft_64_stage_1_0_t1054 * 32 +: 32] = FSM_fft_64_stage_1_0_t1040 - FSM_fft_64_stage_1_0_t1046;
    FSM_fft_64_stage_1_0_t1056 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010000;
    FSM_fft_64_stage_1_0_t1057 = FSM_fft_64_stage_1_0_t1056[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1058 = FSM_fft_64_stage_1_0_t1057[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1059 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010000;
    FSM_fft_64_stage_1_0_t1060 = FSM_fft_64_stage_1_0_t1059[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1061 = FSM_fft_64_stage_1_0_t1060[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1062 = i_data_in_imag[FSM_fft_64_stage_1_0_t1061 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1063 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010000;
    FSM_fft_64_stage_1_0_t1064 = FSM_fft_64_stage_1_0_t1063[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1065 = FSM_fft_64_stage_1_0_t1064 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1066 = FSM_fft_64_stage_1_0_t1065[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1067 = FSM_fft_64_stage_1_0_t1066[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1068 = i_data_in_imag[FSM_fft_64_stage_1_0_t1067 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1069 = FSM_fft_64_stage_1_0_t1062 + FSM_fft_64_stage_1_0_t1068;
    FSM_fft_64_stage_1_0_t1070 = FSM_fft_64_stage_1_0_t1069[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1071 = FSM_fft_64_stage_1_0_t1055;
    FSM_fft_64_stage_1_0_t1071[FSM_fft_64_stage_1_0_t1058 * 32 +: 32] = FSM_fft_64_stage_1_0_t1070;
    FSM_fft_64_stage_1_0_t1072 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010000;
    FSM_fft_64_stage_1_0_t1073 = FSM_fft_64_stage_1_0_t1072[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1074 = FSM_fft_64_stage_1_0_t1073 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1075 = FSM_fft_64_stage_1_0_t1074[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1076 = FSM_fft_64_stage_1_0_t1075[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1077 = FSM_fft_64_stage_1_0_t1071;
    FSM_fft_64_stage_1_0_t1077[FSM_fft_64_stage_1_0_t1076 * 32 +: 32] = FSM_fft_64_stage_1_0_t1062 - FSM_fft_64_stage_1_0_t1068;
    FSM_fft_64_stage_1_0_t1078 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010001;
    FSM_fft_64_stage_1_0_t1079 = FSM_fft_64_stage_1_0_t1078[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1080 = FSM_fft_64_stage_1_0_t1079[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1081 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010001;
    FSM_fft_64_stage_1_0_t1082 = FSM_fft_64_stage_1_0_t1081[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1083 = FSM_fft_64_stage_1_0_t1082[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1084 = i_data_in_imag[FSM_fft_64_stage_1_0_t1083 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1085 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010001;
    FSM_fft_64_stage_1_0_t1086 = FSM_fft_64_stage_1_0_t1085[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1087 = FSM_fft_64_stage_1_0_t1086 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1088 = FSM_fft_64_stage_1_0_t1087[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1089 = FSM_fft_64_stage_1_0_t1088[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1090 = i_data_in_imag[FSM_fft_64_stage_1_0_t1089 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1091 = FSM_fft_64_stage_1_0_t1084 + FSM_fft_64_stage_1_0_t1090;
    FSM_fft_64_stage_1_0_t1092 = FSM_fft_64_stage_1_0_t1091[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1093 = FSM_fft_64_stage_1_0_t1077;
    FSM_fft_64_stage_1_0_t1093[FSM_fft_64_stage_1_0_t1080 * 32 +: 32] = FSM_fft_64_stage_1_0_t1092;
    FSM_fft_64_stage_1_0_t1094 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010001;
    FSM_fft_64_stage_1_0_t1095 = FSM_fft_64_stage_1_0_t1094[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1096 = FSM_fft_64_stage_1_0_t1095 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1097 = FSM_fft_64_stage_1_0_t1096[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1098 = FSM_fft_64_stage_1_0_t1097[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1099 = FSM_fft_64_stage_1_0_t1093;
    FSM_fft_64_stage_1_0_t1099[FSM_fft_64_stage_1_0_t1098 * 32 +: 32] = FSM_fft_64_stage_1_0_t1084 - FSM_fft_64_stage_1_0_t1090;
    FSM_fft_64_stage_1_0_t1100 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010010;
    FSM_fft_64_stage_1_0_t1101 = FSM_fft_64_stage_1_0_t1100[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1102 = FSM_fft_64_stage_1_0_t1101[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1103 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010010;
    FSM_fft_64_stage_1_0_t1104 = FSM_fft_64_stage_1_0_t1103[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1105 = FSM_fft_64_stage_1_0_t1104[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1106 = i_data_in_imag[FSM_fft_64_stage_1_0_t1105 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1107 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010010;
    FSM_fft_64_stage_1_0_t1108 = FSM_fft_64_stage_1_0_t1107[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1109 = FSM_fft_64_stage_1_0_t1108 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1110 = FSM_fft_64_stage_1_0_t1109[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1111 = FSM_fft_64_stage_1_0_t1110[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1112 = i_data_in_imag[FSM_fft_64_stage_1_0_t1111 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1113 = FSM_fft_64_stage_1_0_t1106 + FSM_fft_64_stage_1_0_t1112;
    FSM_fft_64_stage_1_0_t1114 = FSM_fft_64_stage_1_0_t1113[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1115 = FSM_fft_64_stage_1_0_t1099;
    FSM_fft_64_stage_1_0_t1115[FSM_fft_64_stage_1_0_t1102 * 32 +: 32] = FSM_fft_64_stage_1_0_t1114;
    FSM_fft_64_stage_1_0_t1116 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010010;
    FSM_fft_64_stage_1_0_t1117 = FSM_fft_64_stage_1_0_t1116[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1118 = FSM_fft_64_stage_1_0_t1117 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1119 = FSM_fft_64_stage_1_0_t1118[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1120 = FSM_fft_64_stage_1_0_t1119[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1121 = FSM_fft_64_stage_1_0_t1115;
    FSM_fft_64_stage_1_0_t1121[FSM_fft_64_stage_1_0_t1120 * 32 +: 32] = FSM_fft_64_stage_1_0_t1106 - FSM_fft_64_stage_1_0_t1112;
    FSM_fft_64_stage_1_0_t1122 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010011;
    FSM_fft_64_stage_1_0_t1123 = FSM_fft_64_stage_1_0_t1122[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1124 = FSM_fft_64_stage_1_0_t1123[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1125 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010011;
    FSM_fft_64_stage_1_0_t1126 = FSM_fft_64_stage_1_0_t1125[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1127 = FSM_fft_64_stage_1_0_t1126[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1128 = i_data_in_imag[FSM_fft_64_stage_1_0_t1127 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1129 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010011;
    FSM_fft_64_stage_1_0_t1130 = FSM_fft_64_stage_1_0_t1129[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1131 = FSM_fft_64_stage_1_0_t1130 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1132 = FSM_fft_64_stage_1_0_t1131[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1133 = FSM_fft_64_stage_1_0_t1132[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1134 = i_data_in_imag[FSM_fft_64_stage_1_0_t1133 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1135 = FSM_fft_64_stage_1_0_t1128 + FSM_fft_64_stage_1_0_t1134;
    FSM_fft_64_stage_1_0_t1136 = FSM_fft_64_stage_1_0_t1135[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1137 = FSM_fft_64_stage_1_0_t1121;
    FSM_fft_64_stage_1_0_t1137[FSM_fft_64_stage_1_0_t1124 * 32 +: 32] = FSM_fft_64_stage_1_0_t1136;
    FSM_fft_64_stage_1_0_t1138 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010011;
    FSM_fft_64_stage_1_0_t1139 = FSM_fft_64_stage_1_0_t1138[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1140 = FSM_fft_64_stage_1_0_t1139 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1141 = FSM_fft_64_stage_1_0_t1140[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1142 = FSM_fft_64_stage_1_0_t1141[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1143 = FSM_fft_64_stage_1_0_t1137;
    FSM_fft_64_stage_1_0_t1143[FSM_fft_64_stage_1_0_t1142 * 32 +: 32] = FSM_fft_64_stage_1_0_t1128 - FSM_fft_64_stage_1_0_t1134;
    FSM_fft_64_stage_1_0_t1144 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010100;
    FSM_fft_64_stage_1_0_t1145 = FSM_fft_64_stage_1_0_t1144[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1146 = FSM_fft_64_stage_1_0_t1145[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1147 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010100;
    FSM_fft_64_stage_1_0_t1148 = FSM_fft_64_stage_1_0_t1147[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1149 = FSM_fft_64_stage_1_0_t1148[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1150 = i_data_in_imag[FSM_fft_64_stage_1_0_t1149 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1151 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010100;
    FSM_fft_64_stage_1_0_t1152 = FSM_fft_64_stage_1_0_t1151[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1153 = FSM_fft_64_stage_1_0_t1152 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1154 = FSM_fft_64_stage_1_0_t1153[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1155 = FSM_fft_64_stage_1_0_t1154[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1156 = i_data_in_imag[FSM_fft_64_stage_1_0_t1155 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1157 = FSM_fft_64_stage_1_0_t1150 + FSM_fft_64_stage_1_0_t1156;
    FSM_fft_64_stage_1_0_t1158 = FSM_fft_64_stage_1_0_t1157[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1159 = FSM_fft_64_stage_1_0_t1143;
    FSM_fft_64_stage_1_0_t1159[FSM_fft_64_stage_1_0_t1146 * 32 +: 32] = FSM_fft_64_stage_1_0_t1158;
    FSM_fft_64_stage_1_0_t1160 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010100;
    FSM_fft_64_stage_1_0_t1161 = FSM_fft_64_stage_1_0_t1160[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1162 = FSM_fft_64_stage_1_0_t1161 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1163 = FSM_fft_64_stage_1_0_t1162[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1164 = FSM_fft_64_stage_1_0_t1163[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1165 = FSM_fft_64_stage_1_0_t1159;
    FSM_fft_64_stage_1_0_t1165[FSM_fft_64_stage_1_0_t1164 * 32 +: 32] = FSM_fft_64_stage_1_0_t1150 - FSM_fft_64_stage_1_0_t1156;
    FSM_fft_64_stage_1_0_t1166 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010101;
    FSM_fft_64_stage_1_0_t1167 = FSM_fft_64_stage_1_0_t1166[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1168 = FSM_fft_64_stage_1_0_t1167[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1169 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010101;
    FSM_fft_64_stage_1_0_t1170 = FSM_fft_64_stage_1_0_t1169[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1171 = FSM_fft_64_stage_1_0_t1170[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1172 = i_data_in_imag[FSM_fft_64_stage_1_0_t1171 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1173 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010101;
    FSM_fft_64_stage_1_0_t1174 = FSM_fft_64_stage_1_0_t1173[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1175 = FSM_fft_64_stage_1_0_t1174 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1176 = FSM_fft_64_stage_1_0_t1175[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1177 = FSM_fft_64_stage_1_0_t1176[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1178 = i_data_in_imag[FSM_fft_64_stage_1_0_t1177 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1179 = FSM_fft_64_stage_1_0_t1172 + FSM_fft_64_stage_1_0_t1178;
    FSM_fft_64_stage_1_0_t1180 = FSM_fft_64_stage_1_0_t1179[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1181 = FSM_fft_64_stage_1_0_t1165;
    FSM_fft_64_stage_1_0_t1181[FSM_fft_64_stage_1_0_t1168 * 32 +: 32] = FSM_fft_64_stage_1_0_t1180;
    FSM_fft_64_stage_1_0_t1182 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010101;
    FSM_fft_64_stage_1_0_t1183 = FSM_fft_64_stage_1_0_t1182[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1184 = FSM_fft_64_stage_1_0_t1183 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1185 = FSM_fft_64_stage_1_0_t1184[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1186 = FSM_fft_64_stage_1_0_t1185[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1187 = FSM_fft_64_stage_1_0_t1181;
    FSM_fft_64_stage_1_0_t1187[FSM_fft_64_stage_1_0_t1186 * 32 +: 32] = FSM_fft_64_stage_1_0_t1172 - FSM_fft_64_stage_1_0_t1178;
    FSM_fft_64_stage_1_0_t1188 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010110;
    FSM_fft_64_stage_1_0_t1189 = FSM_fft_64_stage_1_0_t1188[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1190 = FSM_fft_64_stage_1_0_t1189[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1191 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010110;
    FSM_fft_64_stage_1_0_t1192 = FSM_fft_64_stage_1_0_t1191[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1193 = FSM_fft_64_stage_1_0_t1192[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1194 = i_data_in_imag[FSM_fft_64_stage_1_0_t1193 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1195 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010110;
    FSM_fft_64_stage_1_0_t1196 = FSM_fft_64_stage_1_0_t1195[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1197 = FSM_fft_64_stage_1_0_t1196 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1198 = FSM_fft_64_stage_1_0_t1197[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1199 = FSM_fft_64_stage_1_0_t1198[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1200 = i_data_in_imag[FSM_fft_64_stage_1_0_t1199 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1201 = FSM_fft_64_stage_1_0_t1194 + FSM_fft_64_stage_1_0_t1200;
    FSM_fft_64_stage_1_0_t1202 = FSM_fft_64_stage_1_0_t1201[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1203 = FSM_fft_64_stage_1_0_t1187;
    FSM_fft_64_stage_1_0_t1203[FSM_fft_64_stage_1_0_t1190 * 32 +: 32] = FSM_fft_64_stage_1_0_t1202;
    FSM_fft_64_stage_1_0_t1204 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010110;
    FSM_fft_64_stage_1_0_t1205 = FSM_fft_64_stage_1_0_t1204[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1206 = FSM_fft_64_stage_1_0_t1205 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1207 = FSM_fft_64_stage_1_0_t1206[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1208 = FSM_fft_64_stage_1_0_t1207[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1209 = FSM_fft_64_stage_1_0_t1203;
    FSM_fft_64_stage_1_0_t1209[FSM_fft_64_stage_1_0_t1208 * 32 +: 32] = FSM_fft_64_stage_1_0_t1194 - FSM_fft_64_stage_1_0_t1200;
    FSM_fft_64_stage_1_0_t1210 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010111;
    FSM_fft_64_stage_1_0_t1211 = FSM_fft_64_stage_1_0_t1210[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1212 = FSM_fft_64_stage_1_0_t1211[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1213 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010111;
    FSM_fft_64_stage_1_0_t1214 = FSM_fft_64_stage_1_0_t1213[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1215 = FSM_fft_64_stage_1_0_t1214[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1216 = i_data_in_imag[FSM_fft_64_stage_1_0_t1215 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1217 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010111;
    FSM_fft_64_stage_1_0_t1218 = FSM_fft_64_stage_1_0_t1217[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1219 = FSM_fft_64_stage_1_0_t1218 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1220 = FSM_fft_64_stage_1_0_t1219[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1221 = FSM_fft_64_stage_1_0_t1220[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1222 = i_data_in_imag[FSM_fft_64_stage_1_0_t1221 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1223 = FSM_fft_64_stage_1_0_t1216 + FSM_fft_64_stage_1_0_t1222;
    FSM_fft_64_stage_1_0_t1224 = FSM_fft_64_stage_1_0_t1223[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1225 = FSM_fft_64_stage_1_0_t1209;
    FSM_fft_64_stage_1_0_t1225[FSM_fft_64_stage_1_0_t1212 * 32 +: 32] = FSM_fft_64_stage_1_0_t1224;
    FSM_fft_64_stage_1_0_t1226 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010111;
    FSM_fft_64_stage_1_0_t1227 = FSM_fft_64_stage_1_0_t1226[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1228 = FSM_fft_64_stage_1_0_t1227 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1229 = FSM_fft_64_stage_1_0_t1228[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1230 = FSM_fft_64_stage_1_0_t1229[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1231 = FSM_fft_64_stage_1_0_t1225;
    FSM_fft_64_stage_1_0_t1231[FSM_fft_64_stage_1_0_t1230 * 32 +: 32] = FSM_fft_64_stage_1_0_t1216 - FSM_fft_64_stage_1_0_t1222;
    FSM_fft_64_stage_1_0_t1232 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011000;
    FSM_fft_64_stage_1_0_t1233 = FSM_fft_64_stage_1_0_t1232[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1234 = FSM_fft_64_stage_1_0_t1233[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1235 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011000;
    FSM_fft_64_stage_1_0_t1236 = FSM_fft_64_stage_1_0_t1235[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1237 = FSM_fft_64_stage_1_0_t1236[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1238 = i_data_in_imag[FSM_fft_64_stage_1_0_t1237 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1239 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011000;
    FSM_fft_64_stage_1_0_t1240 = FSM_fft_64_stage_1_0_t1239[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1241 = FSM_fft_64_stage_1_0_t1240 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1242 = FSM_fft_64_stage_1_0_t1241[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1243 = FSM_fft_64_stage_1_0_t1242[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1244 = i_data_in_imag[FSM_fft_64_stage_1_0_t1243 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1245 = FSM_fft_64_stage_1_0_t1238 + FSM_fft_64_stage_1_0_t1244;
    FSM_fft_64_stage_1_0_t1246 = FSM_fft_64_stage_1_0_t1245[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1247 = FSM_fft_64_stage_1_0_t1231;
    FSM_fft_64_stage_1_0_t1247[FSM_fft_64_stage_1_0_t1234 * 32 +: 32] = FSM_fft_64_stage_1_0_t1246;
    FSM_fft_64_stage_1_0_t1248 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011000;
    FSM_fft_64_stage_1_0_t1249 = FSM_fft_64_stage_1_0_t1248[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1250 = FSM_fft_64_stage_1_0_t1249 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1251 = FSM_fft_64_stage_1_0_t1250[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1252 = FSM_fft_64_stage_1_0_t1251[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1253 = FSM_fft_64_stage_1_0_t1247;
    FSM_fft_64_stage_1_0_t1253[FSM_fft_64_stage_1_0_t1252 * 32 +: 32] = FSM_fft_64_stage_1_0_t1238 - FSM_fft_64_stage_1_0_t1244;
    FSM_fft_64_stage_1_0_t1254 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011001;
    FSM_fft_64_stage_1_0_t1255 = FSM_fft_64_stage_1_0_t1254[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1256 = FSM_fft_64_stage_1_0_t1255[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1257 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011001;
    FSM_fft_64_stage_1_0_t1258 = FSM_fft_64_stage_1_0_t1257[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1259 = FSM_fft_64_stage_1_0_t1258[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1260 = i_data_in_imag[FSM_fft_64_stage_1_0_t1259 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1261 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011001;
    FSM_fft_64_stage_1_0_t1262 = FSM_fft_64_stage_1_0_t1261[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1263 = FSM_fft_64_stage_1_0_t1262 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1264 = FSM_fft_64_stage_1_0_t1263[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1265 = FSM_fft_64_stage_1_0_t1264[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1266 = i_data_in_imag[FSM_fft_64_stage_1_0_t1265 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1267 = FSM_fft_64_stage_1_0_t1260 + FSM_fft_64_stage_1_0_t1266;
    FSM_fft_64_stage_1_0_t1268 = FSM_fft_64_stage_1_0_t1267[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1269 = FSM_fft_64_stage_1_0_t1253;
    FSM_fft_64_stage_1_0_t1269[FSM_fft_64_stage_1_0_t1256 * 32 +: 32] = FSM_fft_64_stage_1_0_t1268;
    FSM_fft_64_stage_1_0_t1270 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011001;
    FSM_fft_64_stage_1_0_t1271 = FSM_fft_64_stage_1_0_t1270[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1272 = FSM_fft_64_stage_1_0_t1271 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1273 = FSM_fft_64_stage_1_0_t1272[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1274 = FSM_fft_64_stage_1_0_t1273[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1275 = FSM_fft_64_stage_1_0_t1269;
    FSM_fft_64_stage_1_0_t1275[FSM_fft_64_stage_1_0_t1274 * 32 +: 32] = FSM_fft_64_stage_1_0_t1260 - FSM_fft_64_stage_1_0_t1266;
    FSM_fft_64_stage_1_0_t1276 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011010;
    FSM_fft_64_stage_1_0_t1277 = FSM_fft_64_stage_1_0_t1276[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1278 = FSM_fft_64_stage_1_0_t1277[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1279 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011010;
    FSM_fft_64_stage_1_0_t1280 = FSM_fft_64_stage_1_0_t1279[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1281 = FSM_fft_64_stage_1_0_t1280[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1282 = i_data_in_imag[FSM_fft_64_stage_1_0_t1281 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1283 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011010;
    FSM_fft_64_stage_1_0_t1284 = FSM_fft_64_stage_1_0_t1283[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1285 = FSM_fft_64_stage_1_0_t1284 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1286 = FSM_fft_64_stage_1_0_t1285[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1287 = FSM_fft_64_stage_1_0_t1286[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1288 = i_data_in_imag[FSM_fft_64_stage_1_0_t1287 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1289 = FSM_fft_64_stage_1_0_t1282 + FSM_fft_64_stage_1_0_t1288;
    FSM_fft_64_stage_1_0_t1290 = FSM_fft_64_stage_1_0_t1289[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1291 = FSM_fft_64_stage_1_0_t1275;
    FSM_fft_64_stage_1_0_t1291[FSM_fft_64_stage_1_0_t1278 * 32 +: 32] = FSM_fft_64_stage_1_0_t1290;
    FSM_fft_64_stage_1_0_t1292 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011010;
    FSM_fft_64_stage_1_0_t1293 = FSM_fft_64_stage_1_0_t1292[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1294 = FSM_fft_64_stage_1_0_t1293 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1295 = FSM_fft_64_stage_1_0_t1294[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1296 = FSM_fft_64_stage_1_0_t1295[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1297 = FSM_fft_64_stage_1_0_t1291;
    FSM_fft_64_stage_1_0_t1297[FSM_fft_64_stage_1_0_t1296 * 32 +: 32] = FSM_fft_64_stage_1_0_t1282 - FSM_fft_64_stage_1_0_t1288;
    FSM_fft_64_stage_1_0_t1298 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011011;
    FSM_fft_64_stage_1_0_t1299 = FSM_fft_64_stage_1_0_t1298[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1300 = FSM_fft_64_stage_1_0_t1299[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1301 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011011;
    FSM_fft_64_stage_1_0_t1302 = FSM_fft_64_stage_1_0_t1301[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1303 = FSM_fft_64_stage_1_0_t1302[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1304 = i_data_in_imag[FSM_fft_64_stage_1_0_t1303 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1305 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011011;
    FSM_fft_64_stage_1_0_t1306 = FSM_fft_64_stage_1_0_t1305[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1307 = FSM_fft_64_stage_1_0_t1306 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1308 = FSM_fft_64_stage_1_0_t1307[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1309 = FSM_fft_64_stage_1_0_t1308[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1310 = i_data_in_imag[FSM_fft_64_stage_1_0_t1309 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1311 = FSM_fft_64_stage_1_0_t1304 + FSM_fft_64_stage_1_0_t1310;
    FSM_fft_64_stage_1_0_t1312 = FSM_fft_64_stage_1_0_t1311[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1313 = FSM_fft_64_stage_1_0_t1297;
    FSM_fft_64_stage_1_0_t1313[FSM_fft_64_stage_1_0_t1300 * 32 +: 32] = FSM_fft_64_stage_1_0_t1312;
    FSM_fft_64_stage_1_0_t1314 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011011;
    FSM_fft_64_stage_1_0_t1315 = FSM_fft_64_stage_1_0_t1314[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1316 = FSM_fft_64_stage_1_0_t1315 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1317 = FSM_fft_64_stage_1_0_t1316[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1318 = FSM_fft_64_stage_1_0_t1317[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1319 = FSM_fft_64_stage_1_0_t1313;
    FSM_fft_64_stage_1_0_t1319[FSM_fft_64_stage_1_0_t1318 * 32 +: 32] = FSM_fft_64_stage_1_0_t1304 - FSM_fft_64_stage_1_0_t1310;
    FSM_fft_64_stage_1_0_t1320 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011100;
    FSM_fft_64_stage_1_0_t1321 = FSM_fft_64_stage_1_0_t1320[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1322 = FSM_fft_64_stage_1_0_t1321[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1323 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011100;
    FSM_fft_64_stage_1_0_t1324 = FSM_fft_64_stage_1_0_t1323[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1325 = FSM_fft_64_stage_1_0_t1324[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1326 = i_data_in_imag[FSM_fft_64_stage_1_0_t1325 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1327 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011100;
    FSM_fft_64_stage_1_0_t1328 = FSM_fft_64_stage_1_0_t1327[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1329 = FSM_fft_64_stage_1_0_t1328 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1330 = FSM_fft_64_stage_1_0_t1329[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1331 = FSM_fft_64_stage_1_0_t1330[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1332 = i_data_in_imag[FSM_fft_64_stage_1_0_t1331 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1333 = FSM_fft_64_stage_1_0_t1326 + FSM_fft_64_stage_1_0_t1332;
    FSM_fft_64_stage_1_0_t1334 = FSM_fft_64_stage_1_0_t1333[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1335 = FSM_fft_64_stage_1_0_t1319;
    FSM_fft_64_stage_1_0_t1335[FSM_fft_64_stage_1_0_t1322 * 32 +: 32] = FSM_fft_64_stage_1_0_t1334;
    FSM_fft_64_stage_1_0_t1336 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011100;
    FSM_fft_64_stage_1_0_t1337 = FSM_fft_64_stage_1_0_t1336[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1338 = FSM_fft_64_stage_1_0_t1337 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1339 = FSM_fft_64_stage_1_0_t1338[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1340 = FSM_fft_64_stage_1_0_t1339[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1341 = FSM_fft_64_stage_1_0_t1335;
    FSM_fft_64_stage_1_0_t1341[FSM_fft_64_stage_1_0_t1340 * 32 +: 32] = FSM_fft_64_stage_1_0_t1326 - FSM_fft_64_stage_1_0_t1332;
    FSM_fft_64_stage_1_0_t1342 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011101;
    FSM_fft_64_stage_1_0_t1343 = FSM_fft_64_stage_1_0_t1342[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1344 = FSM_fft_64_stage_1_0_t1343[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1345 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011101;
    FSM_fft_64_stage_1_0_t1346 = FSM_fft_64_stage_1_0_t1345[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1347 = FSM_fft_64_stage_1_0_t1346[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1348 = i_data_in_imag[FSM_fft_64_stage_1_0_t1347 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1349 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011101;
    FSM_fft_64_stage_1_0_t1350 = FSM_fft_64_stage_1_0_t1349[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1351 = FSM_fft_64_stage_1_0_t1350 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1352 = FSM_fft_64_stage_1_0_t1351[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1353 = FSM_fft_64_stage_1_0_t1352[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1354 = i_data_in_imag[FSM_fft_64_stage_1_0_t1353 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1355 = FSM_fft_64_stage_1_0_t1348 + FSM_fft_64_stage_1_0_t1354;
    FSM_fft_64_stage_1_0_t1356 = FSM_fft_64_stage_1_0_t1355[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1357 = FSM_fft_64_stage_1_0_t1341;
    FSM_fft_64_stage_1_0_t1357[FSM_fft_64_stage_1_0_t1344 * 32 +: 32] = FSM_fft_64_stage_1_0_t1356;
    FSM_fft_64_stage_1_0_t1358 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011101;
    FSM_fft_64_stage_1_0_t1359 = FSM_fft_64_stage_1_0_t1358[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1360 = FSM_fft_64_stage_1_0_t1359 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1361 = FSM_fft_64_stage_1_0_t1360[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1362 = FSM_fft_64_stage_1_0_t1361[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1363 = FSM_fft_64_stage_1_0_t1357;
    FSM_fft_64_stage_1_0_t1363[FSM_fft_64_stage_1_0_t1362 * 32 +: 32] = FSM_fft_64_stage_1_0_t1348 - FSM_fft_64_stage_1_0_t1354;
    FSM_fft_64_stage_1_0_t1364 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011110;
    FSM_fft_64_stage_1_0_t1365 = FSM_fft_64_stage_1_0_t1364[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1366 = FSM_fft_64_stage_1_0_t1365[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1367 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011110;
    FSM_fft_64_stage_1_0_t1368 = FSM_fft_64_stage_1_0_t1367[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1369 = FSM_fft_64_stage_1_0_t1368[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1370 = i_data_in_imag[FSM_fft_64_stage_1_0_t1369 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1371 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011110;
    FSM_fft_64_stage_1_0_t1372 = FSM_fft_64_stage_1_0_t1371[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1373 = FSM_fft_64_stage_1_0_t1372 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1374 = FSM_fft_64_stage_1_0_t1373[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1375 = FSM_fft_64_stage_1_0_t1374[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1376 = i_data_in_imag[FSM_fft_64_stage_1_0_t1375 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1377 = FSM_fft_64_stage_1_0_t1370 + FSM_fft_64_stage_1_0_t1376;
    FSM_fft_64_stage_1_0_t1378 = FSM_fft_64_stage_1_0_t1377[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1379 = FSM_fft_64_stage_1_0_t1363;
    FSM_fft_64_stage_1_0_t1379[FSM_fft_64_stage_1_0_t1366 * 32 +: 32] = FSM_fft_64_stage_1_0_t1378;
    FSM_fft_64_stage_1_0_t1380 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011110;
    FSM_fft_64_stage_1_0_t1381 = FSM_fft_64_stage_1_0_t1380[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1382 = FSM_fft_64_stage_1_0_t1381 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1383 = FSM_fft_64_stage_1_0_t1382[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1384 = FSM_fft_64_stage_1_0_t1383[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1385 = FSM_fft_64_stage_1_0_t1379;
    FSM_fft_64_stage_1_0_t1385[FSM_fft_64_stage_1_0_t1384 * 32 +: 32] = FSM_fft_64_stage_1_0_t1370 - FSM_fft_64_stage_1_0_t1376;
    FSM_fft_64_stage_1_0_t1386 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011111;
    FSM_fft_64_stage_1_0_t1387 = FSM_fft_64_stage_1_0_t1386[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1388 = FSM_fft_64_stage_1_0_t1387[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1389 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011111;
    FSM_fft_64_stage_1_0_t1390 = FSM_fft_64_stage_1_0_t1389[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1391 = FSM_fft_64_stage_1_0_t1390[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1392 = i_data_in_imag[FSM_fft_64_stage_1_0_t1391 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1393 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011111;
    FSM_fft_64_stage_1_0_t1394 = FSM_fft_64_stage_1_0_t1393[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1395 = FSM_fft_64_stage_1_0_t1394 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1396 = FSM_fft_64_stage_1_0_t1395[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1397 = FSM_fft_64_stage_1_0_t1396[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1398 = i_data_in_imag[FSM_fft_64_stage_1_0_t1397 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1399 = FSM_fft_64_stage_1_0_t1392 + FSM_fft_64_stage_1_0_t1398;
    FSM_fft_64_stage_1_0_t1400 = FSM_fft_64_stage_1_0_t1399[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1401 = FSM_fft_64_stage_1_0_t1385;
    FSM_fft_64_stage_1_0_t1401[FSM_fft_64_stage_1_0_t1388 * 32 +: 32] = FSM_fft_64_stage_1_0_t1400;
    FSM_fft_64_stage_1_0_t1402 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011111;
    FSM_fft_64_stage_1_0_t1403 = FSM_fft_64_stage_1_0_t1402[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1404 = FSM_fft_64_stage_1_0_t1403 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1405 = FSM_fft_64_stage_1_0_t1404[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1406 = FSM_fft_64_stage_1_0_t1405[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1407 = FSM_fft_64_stage_1_0_t1401;
    FSM_fft_64_stage_1_0_t1407[FSM_fft_64_stage_1_0_t1406 * 32 +: 32] = FSM_fft_64_stage_1_0_t1392 - FSM_fft_64_stage_1_0_t1398;
end

always @* begin
    FSM_fft_64_stage_1_0_t0 = 32'b00000000000000000000000000000010 * 32'b0;
    FSM_fft_64_stage_1_0_t1 = FSM_fft_64_stage_1_0_t0[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t2 = FSM_fft_64_stage_1_0_t1[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t3 = 32'b00000000000000000000000000000010 * 32'b0;
    FSM_fft_64_stage_1_0_t4 = FSM_fft_64_stage_1_0_t3[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t5 = FSM_fft_64_stage_1_0_t4[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t6 = i_data_in_real[FSM_fft_64_stage_1_0_t5 * 32 +: 32];
    FSM_fft_64_stage_1_0_t7 = 32'b00000000000000000000000000000010 * 32'b0;
    FSM_fft_64_stage_1_0_t8 = FSM_fft_64_stage_1_0_t7[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t9 = FSM_fft_64_stage_1_0_t8 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t10 = FSM_fft_64_stage_1_0_t9[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t11 = FSM_fft_64_stage_1_0_t10[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t12 = i_data_in_real[FSM_fft_64_stage_1_0_t11 * 32 +: 32];
    FSM_fft_64_stage_1_0_t13 = FSM_fft_64_stage_1_0_t6 + FSM_fft_64_stage_1_0_t12;
    FSM_fft_64_stage_1_0_t14 = FSM_fft_64_stage_1_0_t13[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t15 = 2048'b0;
    FSM_fft_64_stage_1_0_t15[FSM_fft_64_stage_1_0_t2 * 32 +: 32] = FSM_fft_64_stage_1_0_t14;
    FSM_fft_64_stage_1_0_t16 = 32'b00000000000000000000000000000010 * 32'b0;
    FSM_fft_64_stage_1_0_t17 = FSM_fft_64_stage_1_0_t16[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t18 = FSM_fft_64_stage_1_0_t17 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t19 = FSM_fft_64_stage_1_0_t18[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t20 = FSM_fft_64_stage_1_0_t19[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t21 = FSM_fft_64_stage_1_0_t15;
    FSM_fft_64_stage_1_0_t21[FSM_fft_64_stage_1_0_t20 * 32 +: 32] = FSM_fft_64_stage_1_0_t6 - FSM_fft_64_stage_1_0_t12;
    FSM_fft_64_stage_1_0_t22 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t23 = FSM_fft_64_stage_1_0_t22[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t24 = FSM_fft_64_stage_1_0_t23[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t25 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t26 = FSM_fft_64_stage_1_0_t25[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t27 = FSM_fft_64_stage_1_0_t26[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t28 = i_data_in_real[FSM_fft_64_stage_1_0_t27 * 32 +: 32];
    FSM_fft_64_stage_1_0_t29 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t30 = FSM_fft_64_stage_1_0_t29[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t31 = FSM_fft_64_stage_1_0_t30 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t32 = FSM_fft_64_stage_1_0_t31[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t33 = FSM_fft_64_stage_1_0_t32[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t34 = i_data_in_real[FSM_fft_64_stage_1_0_t33 * 32 +: 32];
    FSM_fft_64_stage_1_0_t35 = FSM_fft_64_stage_1_0_t28 + FSM_fft_64_stage_1_0_t34;
    FSM_fft_64_stage_1_0_t36 = FSM_fft_64_stage_1_0_t35[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t37 = FSM_fft_64_stage_1_0_t21;
    FSM_fft_64_stage_1_0_t37[FSM_fft_64_stage_1_0_t24 * 32 +: 32] = FSM_fft_64_stage_1_0_t36;
    FSM_fft_64_stage_1_0_t38 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t39 = FSM_fft_64_stage_1_0_t38[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t40 = FSM_fft_64_stage_1_0_t39 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t41 = FSM_fft_64_stage_1_0_t40[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t42 = FSM_fft_64_stage_1_0_t41[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t43 = FSM_fft_64_stage_1_0_t37;
    FSM_fft_64_stage_1_0_t43[FSM_fft_64_stage_1_0_t42 * 32 +: 32] = FSM_fft_64_stage_1_0_t28 - FSM_fft_64_stage_1_0_t34;
    FSM_fft_64_stage_1_0_t44 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_1_0_t45 = FSM_fft_64_stage_1_0_t44[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t46 = FSM_fft_64_stage_1_0_t45[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t47 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_1_0_t48 = FSM_fft_64_stage_1_0_t47[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t49 = FSM_fft_64_stage_1_0_t48[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t50 = i_data_in_real[FSM_fft_64_stage_1_0_t49 * 32 +: 32];
    FSM_fft_64_stage_1_0_t51 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_1_0_t52 = FSM_fft_64_stage_1_0_t51[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t53 = FSM_fft_64_stage_1_0_t52 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t54 = FSM_fft_64_stage_1_0_t53[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t55 = FSM_fft_64_stage_1_0_t54[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t56 = i_data_in_real[FSM_fft_64_stage_1_0_t55 * 32 +: 32];
    FSM_fft_64_stage_1_0_t57 = FSM_fft_64_stage_1_0_t50 + FSM_fft_64_stage_1_0_t56;
    FSM_fft_64_stage_1_0_t58 = FSM_fft_64_stage_1_0_t57[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t59 = FSM_fft_64_stage_1_0_t43;
    FSM_fft_64_stage_1_0_t59[FSM_fft_64_stage_1_0_t46 * 32 +: 32] = FSM_fft_64_stage_1_0_t58;
    FSM_fft_64_stage_1_0_t60 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_1_0_t61 = FSM_fft_64_stage_1_0_t60[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t62 = FSM_fft_64_stage_1_0_t61 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t63 = FSM_fft_64_stage_1_0_t62[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t64 = FSM_fft_64_stage_1_0_t63[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t65 = FSM_fft_64_stage_1_0_t59;
    FSM_fft_64_stage_1_0_t65[FSM_fft_64_stage_1_0_t64 * 32 +: 32] = FSM_fft_64_stage_1_0_t50 - FSM_fft_64_stage_1_0_t56;
    FSM_fft_64_stage_1_0_t66 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_1_0_t67 = FSM_fft_64_stage_1_0_t66[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t68 = FSM_fft_64_stage_1_0_t67[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t69 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_1_0_t70 = FSM_fft_64_stage_1_0_t69[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t71 = FSM_fft_64_stage_1_0_t70[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t72 = i_data_in_real[FSM_fft_64_stage_1_0_t71 * 32 +: 32];
    FSM_fft_64_stage_1_0_t73 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_1_0_t74 = FSM_fft_64_stage_1_0_t73[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t75 = FSM_fft_64_stage_1_0_t74 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t76 = FSM_fft_64_stage_1_0_t75[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t77 = FSM_fft_64_stage_1_0_t76[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t78 = i_data_in_real[FSM_fft_64_stage_1_0_t77 * 32 +: 32];
    FSM_fft_64_stage_1_0_t79 = FSM_fft_64_stage_1_0_t72 + FSM_fft_64_stage_1_0_t78;
    FSM_fft_64_stage_1_0_t80 = FSM_fft_64_stage_1_0_t79[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t81 = FSM_fft_64_stage_1_0_t65;
    FSM_fft_64_stage_1_0_t81[FSM_fft_64_stage_1_0_t68 * 32 +: 32] = FSM_fft_64_stage_1_0_t80;
    FSM_fft_64_stage_1_0_t82 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_1_0_t83 = FSM_fft_64_stage_1_0_t82[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t84 = FSM_fft_64_stage_1_0_t83 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t85 = FSM_fft_64_stage_1_0_t84[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t86 = FSM_fft_64_stage_1_0_t85[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t87 = FSM_fft_64_stage_1_0_t81;
    FSM_fft_64_stage_1_0_t87[FSM_fft_64_stage_1_0_t86 * 32 +: 32] = FSM_fft_64_stage_1_0_t72 - FSM_fft_64_stage_1_0_t78;
    FSM_fft_64_stage_1_0_t88 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000100;
    FSM_fft_64_stage_1_0_t89 = FSM_fft_64_stage_1_0_t88[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t90 = FSM_fft_64_stage_1_0_t89[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t91 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000100;
    FSM_fft_64_stage_1_0_t92 = FSM_fft_64_stage_1_0_t91[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t93 = FSM_fft_64_stage_1_0_t92[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t94 = i_data_in_real[FSM_fft_64_stage_1_0_t93 * 32 +: 32];
    FSM_fft_64_stage_1_0_t95 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000100;
    FSM_fft_64_stage_1_0_t96 = FSM_fft_64_stage_1_0_t95[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t97 = FSM_fft_64_stage_1_0_t96 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t98 = FSM_fft_64_stage_1_0_t97[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t99 = FSM_fft_64_stage_1_0_t98[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t100 = i_data_in_real[FSM_fft_64_stage_1_0_t99 * 32 +: 32];
    FSM_fft_64_stage_1_0_t101 = FSM_fft_64_stage_1_0_t94 + FSM_fft_64_stage_1_0_t100;
    FSM_fft_64_stage_1_0_t102 = FSM_fft_64_stage_1_0_t101[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t103 = FSM_fft_64_stage_1_0_t87;
    FSM_fft_64_stage_1_0_t103[FSM_fft_64_stage_1_0_t90 * 32 +: 32] = FSM_fft_64_stage_1_0_t102;
    FSM_fft_64_stage_1_0_t104 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000100;
    FSM_fft_64_stage_1_0_t105 = FSM_fft_64_stage_1_0_t104[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t106 = FSM_fft_64_stage_1_0_t105 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t107 = FSM_fft_64_stage_1_0_t106[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t108 = FSM_fft_64_stage_1_0_t107[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t109 = FSM_fft_64_stage_1_0_t103;
    FSM_fft_64_stage_1_0_t109[FSM_fft_64_stage_1_0_t108 * 32 +: 32] = FSM_fft_64_stage_1_0_t94 - FSM_fft_64_stage_1_0_t100;
    FSM_fft_64_stage_1_0_t110 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000101;
    FSM_fft_64_stage_1_0_t111 = FSM_fft_64_stage_1_0_t110[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t112 = FSM_fft_64_stage_1_0_t111[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t113 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000101;
    FSM_fft_64_stage_1_0_t114 = FSM_fft_64_stage_1_0_t113[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t115 = FSM_fft_64_stage_1_0_t114[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t116 = i_data_in_real[FSM_fft_64_stage_1_0_t115 * 32 +: 32];
    FSM_fft_64_stage_1_0_t117 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000101;
    FSM_fft_64_stage_1_0_t118 = FSM_fft_64_stage_1_0_t117[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t119 = FSM_fft_64_stage_1_0_t118 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t120 = FSM_fft_64_stage_1_0_t119[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t121 = FSM_fft_64_stage_1_0_t120[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t122 = i_data_in_real[FSM_fft_64_stage_1_0_t121 * 32 +: 32];
    FSM_fft_64_stage_1_0_t123 = FSM_fft_64_stage_1_0_t116 + FSM_fft_64_stage_1_0_t122;
    FSM_fft_64_stage_1_0_t124 = FSM_fft_64_stage_1_0_t123[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t125 = FSM_fft_64_stage_1_0_t109;
    FSM_fft_64_stage_1_0_t125[FSM_fft_64_stage_1_0_t112 * 32 +: 32] = FSM_fft_64_stage_1_0_t124;
    FSM_fft_64_stage_1_0_t126 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000101;
    FSM_fft_64_stage_1_0_t127 = FSM_fft_64_stage_1_0_t126[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t128 = FSM_fft_64_stage_1_0_t127 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t129 = FSM_fft_64_stage_1_0_t128[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t130 = FSM_fft_64_stage_1_0_t129[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t131 = FSM_fft_64_stage_1_0_t125;
    FSM_fft_64_stage_1_0_t131[FSM_fft_64_stage_1_0_t130 * 32 +: 32] = FSM_fft_64_stage_1_0_t116 - FSM_fft_64_stage_1_0_t122;
    FSM_fft_64_stage_1_0_t132 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000110;
    FSM_fft_64_stage_1_0_t133 = FSM_fft_64_stage_1_0_t132[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t134 = FSM_fft_64_stage_1_0_t133[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t135 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000110;
    FSM_fft_64_stage_1_0_t136 = FSM_fft_64_stage_1_0_t135[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t137 = FSM_fft_64_stage_1_0_t136[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t138 = i_data_in_real[FSM_fft_64_stage_1_0_t137 * 32 +: 32];
    FSM_fft_64_stage_1_0_t139 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000110;
    FSM_fft_64_stage_1_0_t140 = FSM_fft_64_stage_1_0_t139[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t141 = FSM_fft_64_stage_1_0_t140 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t142 = FSM_fft_64_stage_1_0_t141[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t143 = FSM_fft_64_stage_1_0_t142[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t144 = i_data_in_real[FSM_fft_64_stage_1_0_t143 * 32 +: 32];
    FSM_fft_64_stage_1_0_t145 = FSM_fft_64_stage_1_0_t138 + FSM_fft_64_stage_1_0_t144;
    FSM_fft_64_stage_1_0_t146 = FSM_fft_64_stage_1_0_t145[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t147 = FSM_fft_64_stage_1_0_t131;
    FSM_fft_64_stage_1_0_t147[FSM_fft_64_stage_1_0_t134 * 32 +: 32] = FSM_fft_64_stage_1_0_t146;
    FSM_fft_64_stage_1_0_t148 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000110;
    FSM_fft_64_stage_1_0_t149 = FSM_fft_64_stage_1_0_t148[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t150 = FSM_fft_64_stage_1_0_t149 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t151 = FSM_fft_64_stage_1_0_t150[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t152 = FSM_fft_64_stage_1_0_t151[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t153 = FSM_fft_64_stage_1_0_t147;
    FSM_fft_64_stage_1_0_t153[FSM_fft_64_stage_1_0_t152 * 32 +: 32] = FSM_fft_64_stage_1_0_t138 - FSM_fft_64_stage_1_0_t144;
    FSM_fft_64_stage_1_0_t154 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000111;
    FSM_fft_64_stage_1_0_t155 = FSM_fft_64_stage_1_0_t154[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t156 = FSM_fft_64_stage_1_0_t155[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t157 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000111;
    FSM_fft_64_stage_1_0_t158 = FSM_fft_64_stage_1_0_t157[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t159 = FSM_fft_64_stage_1_0_t158[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t160 = i_data_in_real[FSM_fft_64_stage_1_0_t159 * 32 +: 32];
    FSM_fft_64_stage_1_0_t161 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000111;
    FSM_fft_64_stage_1_0_t162 = FSM_fft_64_stage_1_0_t161[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t163 = FSM_fft_64_stage_1_0_t162 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t164 = FSM_fft_64_stage_1_0_t163[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t165 = FSM_fft_64_stage_1_0_t164[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t166 = i_data_in_real[FSM_fft_64_stage_1_0_t165 * 32 +: 32];
    FSM_fft_64_stage_1_0_t167 = FSM_fft_64_stage_1_0_t160 + FSM_fft_64_stage_1_0_t166;
    FSM_fft_64_stage_1_0_t168 = FSM_fft_64_stage_1_0_t167[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t169 = FSM_fft_64_stage_1_0_t153;
    FSM_fft_64_stage_1_0_t169[FSM_fft_64_stage_1_0_t156 * 32 +: 32] = FSM_fft_64_stage_1_0_t168;
    FSM_fft_64_stage_1_0_t170 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000111;
    FSM_fft_64_stage_1_0_t171 = FSM_fft_64_stage_1_0_t170[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t172 = FSM_fft_64_stage_1_0_t171 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t173 = FSM_fft_64_stage_1_0_t172[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t174 = FSM_fft_64_stage_1_0_t173[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t175 = FSM_fft_64_stage_1_0_t169;
    FSM_fft_64_stage_1_0_t175[FSM_fft_64_stage_1_0_t174 * 32 +: 32] = FSM_fft_64_stage_1_0_t160 - FSM_fft_64_stage_1_0_t166;
    FSM_fft_64_stage_1_0_t176 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001000;
    FSM_fft_64_stage_1_0_t177 = FSM_fft_64_stage_1_0_t176[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t178 = FSM_fft_64_stage_1_0_t177[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t179 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001000;
    FSM_fft_64_stage_1_0_t180 = FSM_fft_64_stage_1_0_t179[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t181 = FSM_fft_64_stage_1_0_t180[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t182 = i_data_in_real[FSM_fft_64_stage_1_0_t181 * 32 +: 32];
    FSM_fft_64_stage_1_0_t183 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001000;
    FSM_fft_64_stage_1_0_t184 = FSM_fft_64_stage_1_0_t183[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t185 = FSM_fft_64_stage_1_0_t184 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t186 = FSM_fft_64_stage_1_0_t185[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t187 = FSM_fft_64_stage_1_0_t186[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t188 = i_data_in_real[FSM_fft_64_stage_1_0_t187 * 32 +: 32];
    FSM_fft_64_stage_1_0_t189 = FSM_fft_64_stage_1_0_t182 + FSM_fft_64_stage_1_0_t188;
    FSM_fft_64_stage_1_0_t190 = FSM_fft_64_stage_1_0_t189[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t191 = FSM_fft_64_stage_1_0_t175;
    FSM_fft_64_stage_1_0_t191[FSM_fft_64_stage_1_0_t178 * 32 +: 32] = FSM_fft_64_stage_1_0_t190;
    FSM_fft_64_stage_1_0_t192 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001000;
    FSM_fft_64_stage_1_0_t193 = FSM_fft_64_stage_1_0_t192[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t194 = FSM_fft_64_stage_1_0_t193 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t195 = FSM_fft_64_stage_1_0_t194[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t196 = FSM_fft_64_stage_1_0_t195[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t197 = FSM_fft_64_stage_1_0_t191;
    FSM_fft_64_stage_1_0_t197[FSM_fft_64_stage_1_0_t196 * 32 +: 32] = FSM_fft_64_stage_1_0_t182 - FSM_fft_64_stage_1_0_t188;
    FSM_fft_64_stage_1_0_t198 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001001;
    FSM_fft_64_stage_1_0_t199 = FSM_fft_64_stage_1_0_t198[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t200 = FSM_fft_64_stage_1_0_t199[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t201 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001001;
    FSM_fft_64_stage_1_0_t202 = FSM_fft_64_stage_1_0_t201[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t203 = FSM_fft_64_stage_1_0_t202[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t204 = i_data_in_real[FSM_fft_64_stage_1_0_t203 * 32 +: 32];
    FSM_fft_64_stage_1_0_t205 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001001;
    FSM_fft_64_stage_1_0_t206 = FSM_fft_64_stage_1_0_t205[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t207 = FSM_fft_64_stage_1_0_t206 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t208 = FSM_fft_64_stage_1_0_t207[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t209 = FSM_fft_64_stage_1_0_t208[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t210 = i_data_in_real[FSM_fft_64_stage_1_0_t209 * 32 +: 32];
    FSM_fft_64_stage_1_0_t211 = FSM_fft_64_stage_1_0_t204 + FSM_fft_64_stage_1_0_t210;
    FSM_fft_64_stage_1_0_t212 = FSM_fft_64_stage_1_0_t211[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t213 = FSM_fft_64_stage_1_0_t197;
    FSM_fft_64_stage_1_0_t213[FSM_fft_64_stage_1_0_t200 * 32 +: 32] = FSM_fft_64_stage_1_0_t212;
    FSM_fft_64_stage_1_0_t214 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001001;
    FSM_fft_64_stage_1_0_t215 = FSM_fft_64_stage_1_0_t214[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t216 = FSM_fft_64_stage_1_0_t215 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t217 = FSM_fft_64_stage_1_0_t216[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t218 = FSM_fft_64_stage_1_0_t217[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t219 = FSM_fft_64_stage_1_0_t213;
    FSM_fft_64_stage_1_0_t219[FSM_fft_64_stage_1_0_t218 * 32 +: 32] = FSM_fft_64_stage_1_0_t204 - FSM_fft_64_stage_1_0_t210;
    FSM_fft_64_stage_1_0_t220 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001010;
    FSM_fft_64_stage_1_0_t221 = FSM_fft_64_stage_1_0_t220[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t222 = FSM_fft_64_stage_1_0_t221[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t223 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001010;
    FSM_fft_64_stage_1_0_t224 = FSM_fft_64_stage_1_0_t223[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t225 = FSM_fft_64_stage_1_0_t224[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t226 = i_data_in_real[FSM_fft_64_stage_1_0_t225 * 32 +: 32];
    FSM_fft_64_stage_1_0_t227 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001010;
    FSM_fft_64_stage_1_0_t228 = FSM_fft_64_stage_1_0_t227[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t229 = FSM_fft_64_stage_1_0_t228 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t230 = FSM_fft_64_stage_1_0_t229[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t231 = FSM_fft_64_stage_1_0_t230[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t232 = i_data_in_real[FSM_fft_64_stage_1_0_t231 * 32 +: 32];
    FSM_fft_64_stage_1_0_t233 = FSM_fft_64_stage_1_0_t226 + FSM_fft_64_stage_1_0_t232;
    FSM_fft_64_stage_1_0_t234 = FSM_fft_64_stage_1_0_t233[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t235 = FSM_fft_64_stage_1_0_t219;
    FSM_fft_64_stage_1_0_t235[FSM_fft_64_stage_1_0_t222 * 32 +: 32] = FSM_fft_64_stage_1_0_t234;
    FSM_fft_64_stage_1_0_t236 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001010;
    FSM_fft_64_stage_1_0_t237 = FSM_fft_64_stage_1_0_t236[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t238 = FSM_fft_64_stage_1_0_t237 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t239 = FSM_fft_64_stage_1_0_t238[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t240 = FSM_fft_64_stage_1_0_t239[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t241 = FSM_fft_64_stage_1_0_t235;
    FSM_fft_64_stage_1_0_t241[FSM_fft_64_stage_1_0_t240 * 32 +: 32] = FSM_fft_64_stage_1_0_t226 - FSM_fft_64_stage_1_0_t232;
    FSM_fft_64_stage_1_0_t242 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001011;
    FSM_fft_64_stage_1_0_t243 = FSM_fft_64_stage_1_0_t242[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t244 = FSM_fft_64_stage_1_0_t243[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t245 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001011;
    FSM_fft_64_stage_1_0_t246 = FSM_fft_64_stage_1_0_t245[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t247 = FSM_fft_64_stage_1_0_t246[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t248 = i_data_in_real[FSM_fft_64_stage_1_0_t247 * 32 +: 32];
    FSM_fft_64_stage_1_0_t249 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001011;
    FSM_fft_64_stage_1_0_t250 = FSM_fft_64_stage_1_0_t249[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t251 = FSM_fft_64_stage_1_0_t250 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t252 = FSM_fft_64_stage_1_0_t251[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t253 = FSM_fft_64_stage_1_0_t252[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t254 = i_data_in_real[FSM_fft_64_stage_1_0_t253 * 32 +: 32];
    FSM_fft_64_stage_1_0_t255 = FSM_fft_64_stage_1_0_t248 + FSM_fft_64_stage_1_0_t254;
    FSM_fft_64_stage_1_0_t256 = FSM_fft_64_stage_1_0_t255[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t257 = FSM_fft_64_stage_1_0_t241;
    FSM_fft_64_stage_1_0_t257[FSM_fft_64_stage_1_0_t244 * 32 +: 32] = FSM_fft_64_stage_1_0_t256;
    FSM_fft_64_stage_1_0_t258 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001011;
    FSM_fft_64_stage_1_0_t259 = FSM_fft_64_stage_1_0_t258[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t260 = FSM_fft_64_stage_1_0_t259 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t261 = FSM_fft_64_stage_1_0_t260[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t262 = FSM_fft_64_stage_1_0_t261[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t263 = FSM_fft_64_stage_1_0_t257;
    FSM_fft_64_stage_1_0_t263[FSM_fft_64_stage_1_0_t262 * 32 +: 32] = FSM_fft_64_stage_1_0_t248 - FSM_fft_64_stage_1_0_t254;
    FSM_fft_64_stage_1_0_t264 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001100;
    FSM_fft_64_stage_1_0_t265 = FSM_fft_64_stage_1_0_t264[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t266 = FSM_fft_64_stage_1_0_t265[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t267 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001100;
    FSM_fft_64_stage_1_0_t268 = FSM_fft_64_stage_1_0_t267[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t269 = FSM_fft_64_stage_1_0_t268[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t270 = i_data_in_real[FSM_fft_64_stage_1_0_t269 * 32 +: 32];
    FSM_fft_64_stage_1_0_t271 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001100;
    FSM_fft_64_stage_1_0_t272 = FSM_fft_64_stage_1_0_t271[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t273 = FSM_fft_64_stage_1_0_t272 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t274 = FSM_fft_64_stage_1_0_t273[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t275 = FSM_fft_64_stage_1_0_t274[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t276 = i_data_in_real[FSM_fft_64_stage_1_0_t275 * 32 +: 32];
    FSM_fft_64_stage_1_0_t277 = FSM_fft_64_stage_1_0_t270 + FSM_fft_64_stage_1_0_t276;
    FSM_fft_64_stage_1_0_t278 = FSM_fft_64_stage_1_0_t277[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t279 = FSM_fft_64_stage_1_0_t263;
    FSM_fft_64_stage_1_0_t279[FSM_fft_64_stage_1_0_t266 * 32 +: 32] = FSM_fft_64_stage_1_0_t278;
    FSM_fft_64_stage_1_0_t280 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001100;
    FSM_fft_64_stage_1_0_t281 = FSM_fft_64_stage_1_0_t280[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t282 = FSM_fft_64_stage_1_0_t281 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t283 = FSM_fft_64_stage_1_0_t282[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t284 = FSM_fft_64_stage_1_0_t283[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t285 = FSM_fft_64_stage_1_0_t279;
    FSM_fft_64_stage_1_0_t285[FSM_fft_64_stage_1_0_t284 * 32 +: 32] = FSM_fft_64_stage_1_0_t270 - FSM_fft_64_stage_1_0_t276;
    FSM_fft_64_stage_1_0_t286 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001101;
    FSM_fft_64_stage_1_0_t287 = FSM_fft_64_stage_1_0_t286[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t288 = FSM_fft_64_stage_1_0_t287[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t289 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001101;
    FSM_fft_64_stage_1_0_t290 = FSM_fft_64_stage_1_0_t289[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t291 = FSM_fft_64_stage_1_0_t290[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t292 = i_data_in_real[FSM_fft_64_stage_1_0_t291 * 32 +: 32];
    FSM_fft_64_stage_1_0_t293 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001101;
    FSM_fft_64_stage_1_0_t294 = FSM_fft_64_stage_1_0_t293[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t295 = FSM_fft_64_stage_1_0_t294 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t296 = FSM_fft_64_stage_1_0_t295[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t297 = FSM_fft_64_stage_1_0_t296[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t298 = i_data_in_real[FSM_fft_64_stage_1_0_t297 * 32 +: 32];
    FSM_fft_64_stage_1_0_t299 = FSM_fft_64_stage_1_0_t292 + FSM_fft_64_stage_1_0_t298;
    FSM_fft_64_stage_1_0_t300 = FSM_fft_64_stage_1_0_t299[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t301 = FSM_fft_64_stage_1_0_t285;
    FSM_fft_64_stage_1_0_t301[FSM_fft_64_stage_1_0_t288 * 32 +: 32] = FSM_fft_64_stage_1_0_t300;
    FSM_fft_64_stage_1_0_t302 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001101;
    FSM_fft_64_stage_1_0_t303 = FSM_fft_64_stage_1_0_t302[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t304 = FSM_fft_64_stage_1_0_t303 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t305 = FSM_fft_64_stage_1_0_t304[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t306 = FSM_fft_64_stage_1_0_t305[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t307 = FSM_fft_64_stage_1_0_t301;
    FSM_fft_64_stage_1_0_t307[FSM_fft_64_stage_1_0_t306 * 32 +: 32] = FSM_fft_64_stage_1_0_t292 - FSM_fft_64_stage_1_0_t298;
    FSM_fft_64_stage_1_0_t308 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001110;
    FSM_fft_64_stage_1_0_t309 = FSM_fft_64_stage_1_0_t308[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t310 = FSM_fft_64_stage_1_0_t309[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t311 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001110;
    FSM_fft_64_stage_1_0_t312 = FSM_fft_64_stage_1_0_t311[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t313 = FSM_fft_64_stage_1_0_t312[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t314 = i_data_in_real[FSM_fft_64_stage_1_0_t313 * 32 +: 32];
    FSM_fft_64_stage_1_0_t315 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001110;
    FSM_fft_64_stage_1_0_t316 = FSM_fft_64_stage_1_0_t315[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t317 = FSM_fft_64_stage_1_0_t316 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t318 = FSM_fft_64_stage_1_0_t317[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t319 = FSM_fft_64_stage_1_0_t318[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t320 = i_data_in_real[FSM_fft_64_stage_1_0_t319 * 32 +: 32];
    FSM_fft_64_stage_1_0_t321 = FSM_fft_64_stage_1_0_t314 + FSM_fft_64_stage_1_0_t320;
    FSM_fft_64_stage_1_0_t322 = FSM_fft_64_stage_1_0_t321[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t323 = FSM_fft_64_stage_1_0_t307;
    FSM_fft_64_stage_1_0_t323[FSM_fft_64_stage_1_0_t310 * 32 +: 32] = FSM_fft_64_stage_1_0_t322;
    FSM_fft_64_stage_1_0_t324 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001110;
    FSM_fft_64_stage_1_0_t325 = FSM_fft_64_stage_1_0_t324[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t326 = FSM_fft_64_stage_1_0_t325 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t327 = FSM_fft_64_stage_1_0_t326[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t328 = FSM_fft_64_stage_1_0_t327[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t329 = FSM_fft_64_stage_1_0_t323;
    FSM_fft_64_stage_1_0_t329[FSM_fft_64_stage_1_0_t328 * 32 +: 32] = FSM_fft_64_stage_1_0_t314 - FSM_fft_64_stage_1_0_t320;
    FSM_fft_64_stage_1_0_t330 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001111;
    FSM_fft_64_stage_1_0_t331 = FSM_fft_64_stage_1_0_t330[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t332 = FSM_fft_64_stage_1_0_t331[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t333 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001111;
    FSM_fft_64_stage_1_0_t334 = FSM_fft_64_stage_1_0_t333[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t335 = FSM_fft_64_stage_1_0_t334[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t336 = i_data_in_real[FSM_fft_64_stage_1_0_t335 * 32 +: 32];
    FSM_fft_64_stage_1_0_t337 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001111;
    FSM_fft_64_stage_1_0_t338 = FSM_fft_64_stage_1_0_t337[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t339 = FSM_fft_64_stage_1_0_t338 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t340 = FSM_fft_64_stage_1_0_t339[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t341 = FSM_fft_64_stage_1_0_t340[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t342 = i_data_in_real[FSM_fft_64_stage_1_0_t341 * 32 +: 32];
    FSM_fft_64_stage_1_0_t343 = FSM_fft_64_stage_1_0_t336 + FSM_fft_64_stage_1_0_t342;
    FSM_fft_64_stage_1_0_t344 = FSM_fft_64_stage_1_0_t343[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t345 = FSM_fft_64_stage_1_0_t329;
    FSM_fft_64_stage_1_0_t345[FSM_fft_64_stage_1_0_t332 * 32 +: 32] = FSM_fft_64_stage_1_0_t344;
    FSM_fft_64_stage_1_0_t346 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001111;
    FSM_fft_64_stage_1_0_t347 = FSM_fft_64_stage_1_0_t346[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t348 = FSM_fft_64_stage_1_0_t347 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t349 = FSM_fft_64_stage_1_0_t348[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t350 = FSM_fft_64_stage_1_0_t349[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t351 = FSM_fft_64_stage_1_0_t345;
    FSM_fft_64_stage_1_0_t351[FSM_fft_64_stage_1_0_t350 * 32 +: 32] = FSM_fft_64_stage_1_0_t336 - FSM_fft_64_stage_1_0_t342;
    FSM_fft_64_stage_1_0_t352 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010000;
    FSM_fft_64_stage_1_0_t353 = FSM_fft_64_stage_1_0_t352[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t354 = FSM_fft_64_stage_1_0_t353[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t355 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010000;
    FSM_fft_64_stage_1_0_t356 = FSM_fft_64_stage_1_0_t355[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t357 = FSM_fft_64_stage_1_0_t356[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t358 = i_data_in_real[FSM_fft_64_stage_1_0_t357 * 32 +: 32];
    FSM_fft_64_stage_1_0_t359 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010000;
    FSM_fft_64_stage_1_0_t360 = FSM_fft_64_stage_1_0_t359[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t361 = FSM_fft_64_stage_1_0_t360 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t362 = FSM_fft_64_stage_1_0_t361[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t363 = FSM_fft_64_stage_1_0_t362[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t364 = i_data_in_real[FSM_fft_64_stage_1_0_t363 * 32 +: 32];
    FSM_fft_64_stage_1_0_t365 = FSM_fft_64_stage_1_0_t358 + FSM_fft_64_stage_1_0_t364;
    FSM_fft_64_stage_1_0_t366 = FSM_fft_64_stage_1_0_t365[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t367 = FSM_fft_64_stage_1_0_t351;
    FSM_fft_64_stage_1_0_t367[FSM_fft_64_stage_1_0_t354 * 32 +: 32] = FSM_fft_64_stage_1_0_t366;
    FSM_fft_64_stage_1_0_t368 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010000;
    FSM_fft_64_stage_1_0_t369 = FSM_fft_64_stage_1_0_t368[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t370 = FSM_fft_64_stage_1_0_t369 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t371 = FSM_fft_64_stage_1_0_t370[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t372 = FSM_fft_64_stage_1_0_t371[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t373 = FSM_fft_64_stage_1_0_t367;
    FSM_fft_64_stage_1_0_t373[FSM_fft_64_stage_1_0_t372 * 32 +: 32] = FSM_fft_64_stage_1_0_t358 - FSM_fft_64_stage_1_0_t364;
    FSM_fft_64_stage_1_0_t374 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010001;
    FSM_fft_64_stage_1_0_t375 = FSM_fft_64_stage_1_0_t374[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t376 = FSM_fft_64_stage_1_0_t375[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t377 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010001;
    FSM_fft_64_stage_1_0_t378 = FSM_fft_64_stage_1_0_t377[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t379 = FSM_fft_64_stage_1_0_t378[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t380 = i_data_in_real[FSM_fft_64_stage_1_0_t379 * 32 +: 32];
    FSM_fft_64_stage_1_0_t381 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010001;
    FSM_fft_64_stage_1_0_t382 = FSM_fft_64_stage_1_0_t381[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t383 = FSM_fft_64_stage_1_0_t382 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t384 = FSM_fft_64_stage_1_0_t383[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t385 = FSM_fft_64_stage_1_0_t384[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t386 = i_data_in_real[FSM_fft_64_stage_1_0_t385 * 32 +: 32];
    FSM_fft_64_stage_1_0_t387 = FSM_fft_64_stage_1_0_t380 + FSM_fft_64_stage_1_0_t386;
    FSM_fft_64_stage_1_0_t388 = FSM_fft_64_stage_1_0_t387[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t389 = FSM_fft_64_stage_1_0_t373;
    FSM_fft_64_stage_1_0_t389[FSM_fft_64_stage_1_0_t376 * 32 +: 32] = FSM_fft_64_stage_1_0_t388;
    FSM_fft_64_stage_1_0_t390 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010001;
    FSM_fft_64_stage_1_0_t391 = FSM_fft_64_stage_1_0_t390[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t392 = FSM_fft_64_stage_1_0_t391 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t393 = FSM_fft_64_stage_1_0_t392[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t394 = FSM_fft_64_stage_1_0_t393[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t395 = FSM_fft_64_stage_1_0_t389;
    FSM_fft_64_stage_1_0_t395[FSM_fft_64_stage_1_0_t394 * 32 +: 32] = FSM_fft_64_stage_1_0_t380 - FSM_fft_64_stage_1_0_t386;
    FSM_fft_64_stage_1_0_t396 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010010;
    FSM_fft_64_stage_1_0_t397 = FSM_fft_64_stage_1_0_t396[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t398 = FSM_fft_64_stage_1_0_t397[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t399 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010010;
    FSM_fft_64_stage_1_0_t400 = FSM_fft_64_stage_1_0_t399[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t401 = FSM_fft_64_stage_1_0_t400[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t402 = i_data_in_real[FSM_fft_64_stage_1_0_t401 * 32 +: 32];
    FSM_fft_64_stage_1_0_t403 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010010;
    FSM_fft_64_stage_1_0_t404 = FSM_fft_64_stage_1_0_t403[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t405 = FSM_fft_64_stage_1_0_t404 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t406 = FSM_fft_64_stage_1_0_t405[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t407 = FSM_fft_64_stage_1_0_t406[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t408 = i_data_in_real[FSM_fft_64_stage_1_0_t407 * 32 +: 32];
    FSM_fft_64_stage_1_0_t409 = FSM_fft_64_stage_1_0_t402 + FSM_fft_64_stage_1_0_t408;
    FSM_fft_64_stage_1_0_t410 = FSM_fft_64_stage_1_0_t409[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t411 = FSM_fft_64_stage_1_0_t395;
    FSM_fft_64_stage_1_0_t411[FSM_fft_64_stage_1_0_t398 * 32 +: 32] = FSM_fft_64_stage_1_0_t410;
    FSM_fft_64_stage_1_0_t412 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010010;
    FSM_fft_64_stage_1_0_t413 = FSM_fft_64_stage_1_0_t412[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t414 = FSM_fft_64_stage_1_0_t413 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t415 = FSM_fft_64_stage_1_0_t414[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t416 = FSM_fft_64_stage_1_0_t415[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t417 = FSM_fft_64_stage_1_0_t411;
    FSM_fft_64_stage_1_0_t417[FSM_fft_64_stage_1_0_t416 * 32 +: 32] = FSM_fft_64_stage_1_0_t402 - FSM_fft_64_stage_1_0_t408;
    FSM_fft_64_stage_1_0_t418 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010011;
    FSM_fft_64_stage_1_0_t419 = FSM_fft_64_stage_1_0_t418[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t420 = FSM_fft_64_stage_1_0_t419[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t421 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010011;
    FSM_fft_64_stage_1_0_t422 = FSM_fft_64_stage_1_0_t421[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t423 = FSM_fft_64_stage_1_0_t422[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t424 = i_data_in_real[FSM_fft_64_stage_1_0_t423 * 32 +: 32];
    FSM_fft_64_stage_1_0_t425 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010011;
    FSM_fft_64_stage_1_0_t426 = FSM_fft_64_stage_1_0_t425[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t427 = FSM_fft_64_stage_1_0_t426 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t428 = FSM_fft_64_stage_1_0_t427[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t429 = FSM_fft_64_stage_1_0_t428[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t430 = i_data_in_real[FSM_fft_64_stage_1_0_t429 * 32 +: 32];
    FSM_fft_64_stage_1_0_t431 = FSM_fft_64_stage_1_0_t424 + FSM_fft_64_stage_1_0_t430;
    FSM_fft_64_stage_1_0_t432 = FSM_fft_64_stage_1_0_t431[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t433 = FSM_fft_64_stage_1_0_t417;
    FSM_fft_64_stage_1_0_t433[FSM_fft_64_stage_1_0_t420 * 32 +: 32] = FSM_fft_64_stage_1_0_t432;
    FSM_fft_64_stage_1_0_t434 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010011;
    FSM_fft_64_stage_1_0_t435 = FSM_fft_64_stage_1_0_t434[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t436 = FSM_fft_64_stage_1_0_t435 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t437 = FSM_fft_64_stage_1_0_t436[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t438 = FSM_fft_64_stage_1_0_t437[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t439 = FSM_fft_64_stage_1_0_t433;
    FSM_fft_64_stage_1_0_t439[FSM_fft_64_stage_1_0_t438 * 32 +: 32] = FSM_fft_64_stage_1_0_t424 - FSM_fft_64_stage_1_0_t430;
    FSM_fft_64_stage_1_0_t440 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010100;
    FSM_fft_64_stage_1_0_t441 = FSM_fft_64_stage_1_0_t440[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t442 = FSM_fft_64_stage_1_0_t441[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t443 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010100;
    FSM_fft_64_stage_1_0_t444 = FSM_fft_64_stage_1_0_t443[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t445 = FSM_fft_64_stage_1_0_t444[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t446 = i_data_in_real[FSM_fft_64_stage_1_0_t445 * 32 +: 32];
    FSM_fft_64_stage_1_0_t447 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010100;
    FSM_fft_64_stage_1_0_t448 = FSM_fft_64_stage_1_0_t447[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t449 = FSM_fft_64_stage_1_0_t448 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t450 = FSM_fft_64_stage_1_0_t449[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t451 = FSM_fft_64_stage_1_0_t450[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t452 = i_data_in_real[FSM_fft_64_stage_1_0_t451 * 32 +: 32];
    FSM_fft_64_stage_1_0_t453 = FSM_fft_64_stage_1_0_t446 + FSM_fft_64_stage_1_0_t452;
    FSM_fft_64_stage_1_0_t454 = FSM_fft_64_stage_1_0_t453[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t455 = FSM_fft_64_stage_1_0_t439;
    FSM_fft_64_stage_1_0_t455[FSM_fft_64_stage_1_0_t442 * 32 +: 32] = FSM_fft_64_stage_1_0_t454;
    FSM_fft_64_stage_1_0_t456 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010100;
    FSM_fft_64_stage_1_0_t457 = FSM_fft_64_stage_1_0_t456[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t458 = FSM_fft_64_stage_1_0_t457 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t459 = FSM_fft_64_stage_1_0_t458[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t460 = FSM_fft_64_stage_1_0_t459[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t461 = FSM_fft_64_stage_1_0_t455;
    FSM_fft_64_stage_1_0_t461[FSM_fft_64_stage_1_0_t460 * 32 +: 32] = FSM_fft_64_stage_1_0_t446 - FSM_fft_64_stage_1_0_t452;
    FSM_fft_64_stage_1_0_t462 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010101;
    FSM_fft_64_stage_1_0_t463 = FSM_fft_64_stage_1_0_t462[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t464 = FSM_fft_64_stage_1_0_t463[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t465 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010101;
    FSM_fft_64_stage_1_0_t466 = FSM_fft_64_stage_1_0_t465[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t467 = FSM_fft_64_stage_1_0_t466[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t468 = i_data_in_real[FSM_fft_64_stage_1_0_t467 * 32 +: 32];
    FSM_fft_64_stage_1_0_t469 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010101;
    FSM_fft_64_stage_1_0_t470 = FSM_fft_64_stage_1_0_t469[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t471 = FSM_fft_64_stage_1_0_t470 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t472 = FSM_fft_64_stage_1_0_t471[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t473 = FSM_fft_64_stage_1_0_t472[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t474 = i_data_in_real[FSM_fft_64_stage_1_0_t473 * 32 +: 32];
    FSM_fft_64_stage_1_0_t475 = FSM_fft_64_stage_1_0_t468 + FSM_fft_64_stage_1_0_t474;
    FSM_fft_64_stage_1_0_t476 = FSM_fft_64_stage_1_0_t475[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t477 = FSM_fft_64_stage_1_0_t461;
    FSM_fft_64_stage_1_0_t477[FSM_fft_64_stage_1_0_t464 * 32 +: 32] = FSM_fft_64_stage_1_0_t476;
    FSM_fft_64_stage_1_0_t478 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010101;
    FSM_fft_64_stage_1_0_t479 = FSM_fft_64_stage_1_0_t478[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t480 = FSM_fft_64_stage_1_0_t479 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t481 = FSM_fft_64_stage_1_0_t480[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t482 = FSM_fft_64_stage_1_0_t481[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t483 = FSM_fft_64_stage_1_0_t477;
    FSM_fft_64_stage_1_0_t483[FSM_fft_64_stage_1_0_t482 * 32 +: 32] = FSM_fft_64_stage_1_0_t468 - FSM_fft_64_stage_1_0_t474;
    FSM_fft_64_stage_1_0_t484 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010110;
    FSM_fft_64_stage_1_0_t485 = FSM_fft_64_stage_1_0_t484[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t486 = FSM_fft_64_stage_1_0_t485[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t487 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010110;
    FSM_fft_64_stage_1_0_t488 = FSM_fft_64_stage_1_0_t487[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t489 = FSM_fft_64_stage_1_0_t488[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t490 = i_data_in_real[FSM_fft_64_stage_1_0_t489 * 32 +: 32];
    FSM_fft_64_stage_1_0_t491 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010110;
    FSM_fft_64_stage_1_0_t492 = FSM_fft_64_stage_1_0_t491[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t493 = FSM_fft_64_stage_1_0_t492 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t494 = FSM_fft_64_stage_1_0_t493[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t495 = FSM_fft_64_stage_1_0_t494[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t496 = i_data_in_real[FSM_fft_64_stage_1_0_t495 * 32 +: 32];
    FSM_fft_64_stage_1_0_t497 = FSM_fft_64_stage_1_0_t490 + FSM_fft_64_stage_1_0_t496;
    FSM_fft_64_stage_1_0_t498 = FSM_fft_64_stage_1_0_t497[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t499 = FSM_fft_64_stage_1_0_t483;
    FSM_fft_64_stage_1_0_t499[FSM_fft_64_stage_1_0_t486 * 32 +: 32] = FSM_fft_64_stage_1_0_t498;
    FSM_fft_64_stage_1_0_t500 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010110;
    FSM_fft_64_stage_1_0_t501 = FSM_fft_64_stage_1_0_t500[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t502 = FSM_fft_64_stage_1_0_t501 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t503 = FSM_fft_64_stage_1_0_t502[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t504 = FSM_fft_64_stage_1_0_t503[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t505 = FSM_fft_64_stage_1_0_t499;
    FSM_fft_64_stage_1_0_t505[FSM_fft_64_stage_1_0_t504 * 32 +: 32] = FSM_fft_64_stage_1_0_t490 - FSM_fft_64_stage_1_0_t496;
    FSM_fft_64_stage_1_0_t506 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010111;
    FSM_fft_64_stage_1_0_t507 = FSM_fft_64_stage_1_0_t506[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t508 = FSM_fft_64_stage_1_0_t507[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t509 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010111;
    FSM_fft_64_stage_1_0_t510 = FSM_fft_64_stage_1_0_t509[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t511 = FSM_fft_64_stage_1_0_t510[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t512 = i_data_in_real[FSM_fft_64_stage_1_0_t511 * 32 +: 32];
    FSM_fft_64_stage_1_0_t513 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010111;
    FSM_fft_64_stage_1_0_t514 = FSM_fft_64_stage_1_0_t513[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t515 = FSM_fft_64_stage_1_0_t514 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t516 = FSM_fft_64_stage_1_0_t515[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t517 = FSM_fft_64_stage_1_0_t516[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t518 = i_data_in_real[FSM_fft_64_stage_1_0_t517 * 32 +: 32];
    FSM_fft_64_stage_1_0_t519 = FSM_fft_64_stage_1_0_t512 + FSM_fft_64_stage_1_0_t518;
    FSM_fft_64_stage_1_0_t520 = FSM_fft_64_stage_1_0_t519[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t521 = FSM_fft_64_stage_1_0_t505;
    FSM_fft_64_stage_1_0_t521[FSM_fft_64_stage_1_0_t508 * 32 +: 32] = FSM_fft_64_stage_1_0_t520;
    FSM_fft_64_stage_1_0_t522 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010111;
    FSM_fft_64_stage_1_0_t523 = FSM_fft_64_stage_1_0_t522[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t524 = FSM_fft_64_stage_1_0_t523 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t525 = FSM_fft_64_stage_1_0_t524[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t526 = FSM_fft_64_stage_1_0_t525[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t527 = FSM_fft_64_stage_1_0_t521;
    FSM_fft_64_stage_1_0_t527[FSM_fft_64_stage_1_0_t526 * 32 +: 32] = FSM_fft_64_stage_1_0_t512 - FSM_fft_64_stage_1_0_t518;
    FSM_fft_64_stage_1_0_t528 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011000;
    FSM_fft_64_stage_1_0_t529 = FSM_fft_64_stage_1_0_t528[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t530 = FSM_fft_64_stage_1_0_t529[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t531 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011000;
    FSM_fft_64_stage_1_0_t532 = FSM_fft_64_stage_1_0_t531[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t533 = FSM_fft_64_stage_1_0_t532[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t534 = i_data_in_real[FSM_fft_64_stage_1_0_t533 * 32 +: 32];
    FSM_fft_64_stage_1_0_t535 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011000;
    FSM_fft_64_stage_1_0_t536 = FSM_fft_64_stage_1_0_t535[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t537 = FSM_fft_64_stage_1_0_t536 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t538 = FSM_fft_64_stage_1_0_t537[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t539 = FSM_fft_64_stage_1_0_t538[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t540 = i_data_in_real[FSM_fft_64_stage_1_0_t539 * 32 +: 32];
    FSM_fft_64_stage_1_0_t541 = FSM_fft_64_stage_1_0_t534 + FSM_fft_64_stage_1_0_t540;
    FSM_fft_64_stage_1_0_t542 = FSM_fft_64_stage_1_0_t541[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t543 = FSM_fft_64_stage_1_0_t527;
    FSM_fft_64_stage_1_0_t543[FSM_fft_64_stage_1_0_t530 * 32 +: 32] = FSM_fft_64_stage_1_0_t542;
    FSM_fft_64_stage_1_0_t544 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011000;
    FSM_fft_64_stage_1_0_t545 = FSM_fft_64_stage_1_0_t544[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t546 = FSM_fft_64_stage_1_0_t545 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t547 = FSM_fft_64_stage_1_0_t546[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t548 = FSM_fft_64_stage_1_0_t547[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t549 = FSM_fft_64_stage_1_0_t543;
    FSM_fft_64_stage_1_0_t549[FSM_fft_64_stage_1_0_t548 * 32 +: 32] = FSM_fft_64_stage_1_0_t534 - FSM_fft_64_stage_1_0_t540;
    FSM_fft_64_stage_1_0_t550 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011001;
    FSM_fft_64_stage_1_0_t551 = FSM_fft_64_stage_1_0_t550[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t552 = FSM_fft_64_stage_1_0_t551[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t553 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011001;
    FSM_fft_64_stage_1_0_t554 = FSM_fft_64_stage_1_0_t553[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t555 = FSM_fft_64_stage_1_0_t554[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t556 = i_data_in_real[FSM_fft_64_stage_1_0_t555 * 32 +: 32];
    FSM_fft_64_stage_1_0_t557 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011001;
    FSM_fft_64_stage_1_0_t558 = FSM_fft_64_stage_1_0_t557[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t559 = FSM_fft_64_stage_1_0_t558 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t560 = FSM_fft_64_stage_1_0_t559[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t561 = FSM_fft_64_stage_1_0_t560[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t562 = i_data_in_real[FSM_fft_64_stage_1_0_t561 * 32 +: 32];
    FSM_fft_64_stage_1_0_t563 = FSM_fft_64_stage_1_0_t556 + FSM_fft_64_stage_1_0_t562;
    FSM_fft_64_stage_1_0_t564 = FSM_fft_64_stage_1_0_t563[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t565 = FSM_fft_64_stage_1_0_t549;
    FSM_fft_64_stage_1_0_t565[FSM_fft_64_stage_1_0_t552 * 32 +: 32] = FSM_fft_64_stage_1_0_t564;
    FSM_fft_64_stage_1_0_t566 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011001;
    FSM_fft_64_stage_1_0_t567 = FSM_fft_64_stage_1_0_t566[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t568 = FSM_fft_64_stage_1_0_t567 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t569 = FSM_fft_64_stage_1_0_t568[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t570 = FSM_fft_64_stage_1_0_t569[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t571 = FSM_fft_64_stage_1_0_t565;
    FSM_fft_64_stage_1_0_t571[FSM_fft_64_stage_1_0_t570 * 32 +: 32] = FSM_fft_64_stage_1_0_t556 - FSM_fft_64_stage_1_0_t562;
    FSM_fft_64_stage_1_0_t572 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011010;
    FSM_fft_64_stage_1_0_t573 = FSM_fft_64_stage_1_0_t572[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t574 = FSM_fft_64_stage_1_0_t573[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t575 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011010;
    FSM_fft_64_stage_1_0_t576 = FSM_fft_64_stage_1_0_t575[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t577 = FSM_fft_64_stage_1_0_t576[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t578 = i_data_in_real[FSM_fft_64_stage_1_0_t577 * 32 +: 32];
    FSM_fft_64_stage_1_0_t579 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011010;
    FSM_fft_64_stage_1_0_t580 = FSM_fft_64_stage_1_0_t579[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t581 = FSM_fft_64_stage_1_0_t580 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t582 = FSM_fft_64_stage_1_0_t581[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t583 = FSM_fft_64_stage_1_0_t582[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t584 = i_data_in_real[FSM_fft_64_stage_1_0_t583 * 32 +: 32];
    FSM_fft_64_stage_1_0_t585 = FSM_fft_64_stage_1_0_t578 + FSM_fft_64_stage_1_0_t584;
    FSM_fft_64_stage_1_0_t586 = FSM_fft_64_stage_1_0_t585[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t587 = FSM_fft_64_stage_1_0_t571;
    FSM_fft_64_stage_1_0_t587[FSM_fft_64_stage_1_0_t574 * 32 +: 32] = FSM_fft_64_stage_1_0_t586;
    FSM_fft_64_stage_1_0_t588 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011010;
    FSM_fft_64_stage_1_0_t589 = FSM_fft_64_stage_1_0_t588[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t590 = FSM_fft_64_stage_1_0_t589 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t591 = FSM_fft_64_stage_1_0_t590[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t592 = FSM_fft_64_stage_1_0_t591[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t593 = FSM_fft_64_stage_1_0_t587;
    FSM_fft_64_stage_1_0_t593[FSM_fft_64_stage_1_0_t592 * 32 +: 32] = FSM_fft_64_stage_1_0_t578 - FSM_fft_64_stage_1_0_t584;
    FSM_fft_64_stage_1_0_t594 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011011;
    FSM_fft_64_stage_1_0_t595 = FSM_fft_64_stage_1_0_t594[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t596 = FSM_fft_64_stage_1_0_t595[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t597 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011011;
    FSM_fft_64_stage_1_0_t598 = FSM_fft_64_stage_1_0_t597[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t599 = FSM_fft_64_stage_1_0_t598[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t600 = i_data_in_real[FSM_fft_64_stage_1_0_t599 * 32 +: 32];
    FSM_fft_64_stage_1_0_t601 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011011;
    FSM_fft_64_stage_1_0_t602 = FSM_fft_64_stage_1_0_t601[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t603 = FSM_fft_64_stage_1_0_t602 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t604 = FSM_fft_64_stage_1_0_t603[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t605 = FSM_fft_64_stage_1_0_t604[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t606 = i_data_in_real[FSM_fft_64_stage_1_0_t605 * 32 +: 32];
    FSM_fft_64_stage_1_0_t607 = FSM_fft_64_stage_1_0_t600 + FSM_fft_64_stage_1_0_t606;
    FSM_fft_64_stage_1_0_t608 = FSM_fft_64_stage_1_0_t607[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t609 = FSM_fft_64_stage_1_0_t593;
    FSM_fft_64_stage_1_0_t609[FSM_fft_64_stage_1_0_t596 * 32 +: 32] = FSM_fft_64_stage_1_0_t608;
    FSM_fft_64_stage_1_0_t610 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011011;
    FSM_fft_64_stage_1_0_t611 = FSM_fft_64_stage_1_0_t610[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t612 = FSM_fft_64_stage_1_0_t611 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t613 = FSM_fft_64_stage_1_0_t612[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t614 = FSM_fft_64_stage_1_0_t613[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t615 = FSM_fft_64_stage_1_0_t609;
    FSM_fft_64_stage_1_0_t615[FSM_fft_64_stage_1_0_t614 * 32 +: 32] = FSM_fft_64_stage_1_0_t600 - FSM_fft_64_stage_1_0_t606;
    FSM_fft_64_stage_1_0_t616 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011100;
    FSM_fft_64_stage_1_0_t617 = FSM_fft_64_stage_1_0_t616[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t618 = FSM_fft_64_stage_1_0_t617[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t619 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011100;
    FSM_fft_64_stage_1_0_t620 = FSM_fft_64_stage_1_0_t619[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t621 = FSM_fft_64_stage_1_0_t620[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t622 = i_data_in_real[FSM_fft_64_stage_1_0_t621 * 32 +: 32];
    FSM_fft_64_stage_1_0_t623 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011100;
    FSM_fft_64_stage_1_0_t624 = FSM_fft_64_stage_1_0_t623[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t625 = FSM_fft_64_stage_1_0_t624 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t626 = FSM_fft_64_stage_1_0_t625[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t627 = FSM_fft_64_stage_1_0_t626[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t628 = i_data_in_real[FSM_fft_64_stage_1_0_t627 * 32 +: 32];
    FSM_fft_64_stage_1_0_t629 = FSM_fft_64_stage_1_0_t622 + FSM_fft_64_stage_1_0_t628;
    FSM_fft_64_stage_1_0_t630 = FSM_fft_64_stage_1_0_t629[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t631 = FSM_fft_64_stage_1_0_t615;
    FSM_fft_64_stage_1_0_t631[FSM_fft_64_stage_1_0_t618 * 32 +: 32] = FSM_fft_64_stage_1_0_t630;
    FSM_fft_64_stage_1_0_t632 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011100;
    FSM_fft_64_stage_1_0_t633 = FSM_fft_64_stage_1_0_t632[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t634 = FSM_fft_64_stage_1_0_t633 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t635 = FSM_fft_64_stage_1_0_t634[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t636 = FSM_fft_64_stage_1_0_t635[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t637 = FSM_fft_64_stage_1_0_t631;
    FSM_fft_64_stage_1_0_t637[FSM_fft_64_stage_1_0_t636 * 32 +: 32] = FSM_fft_64_stage_1_0_t622 - FSM_fft_64_stage_1_0_t628;
    FSM_fft_64_stage_1_0_t638 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011101;
    FSM_fft_64_stage_1_0_t639 = FSM_fft_64_stage_1_0_t638[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t640 = FSM_fft_64_stage_1_0_t639[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t641 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011101;
    FSM_fft_64_stage_1_0_t642 = FSM_fft_64_stage_1_0_t641[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t643 = FSM_fft_64_stage_1_0_t642[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t644 = i_data_in_real[FSM_fft_64_stage_1_0_t643 * 32 +: 32];
    FSM_fft_64_stage_1_0_t645 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011101;
    FSM_fft_64_stage_1_0_t646 = FSM_fft_64_stage_1_0_t645[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t647 = FSM_fft_64_stage_1_0_t646 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t648 = FSM_fft_64_stage_1_0_t647[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t649 = FSM_fft_64_stage_1_0_t648[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t650 = i_data_in_real[FSM_fft_64_stage_1_0_t649 * 32 +: 32];
    FSM_fft_64_stage_1_0_t651 = FSM_fft_64_stage_1_0_t644 + FSM_fft_64_stage_1_0_t650;
    FSM_fft_64_stage_1_0_t652 = FSM_fft_64_stage_1_0_t651[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t653 = FSM_fft_64_stage_1_0_t637;
    FSM_fft_64_stage_1_0_t653[FSM_fft_64_stage_1_0_t640 * 32 +: 32] = FSM_fft_64_stage_1_0_t652;
    FSM_fft_64_stage_1_0_t654 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011101;
    FSM_fft_64_stage_1_0_t655 = FSM_fft_64_stage_1_0_t654[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t656 = FSM_fft_64_stage_1_0_t655 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t657 = FSM_fft_64_stage_1_0_t656[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t658 = FSM_fft_64_stage_1_0_t657[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t659 = FSM_fft_64_stage_1_0_t653;
    FSM_fft_64_stage_1_0_t659[FSM_fft_64_stage_1_0_t658 * 32 +: 32] = FSM_fft_64_stage_1_0_t644 - FSM_fft_64_stage_1_0_t650;
    FSM_fft_64_stage_1_0_t660 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011110;
    FSM_fft_64_stage_1_0_t661 = FSM_fft_64_stage_1_0_t660[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t662 = FSM_fft_64_stage_1_0_t661[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t663 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011110;
    FSM_fft_64_stage_1_0_t664 = FSM_fft_64_stage_1_0_t663[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t665 = FSM_fft_64_stage_1_0_t664[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t666 = i_data_in_real[FSM_fft_64_stage_1_0_t665 * 32 +: 32];
    FSM_fft_64_stage_1_0_t667 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011110;
    FSM_fft_64_stage_1_0_t668 = FSM_fft_64_stage_1_0_t667[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t669 = FSM_fft_64_stage_1_0_t668 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t670 = FSM_fft_64_stage_1_0_t669[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t671 = FSM_fft_64_stage_1_0_t670[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t672 = i_data_in_real[FSM_fft_64_stage_1_0_t671 * 32 +: 32];
    FSM_fft_64_stage_1_0_t673 = FSM_fft_64_stage_1_0_t666 + FSM_fft_64_stage_1_0_t672;
    FSM_fft_64_stage_1_0_t674 = FSM_fft_64_stage_1_0_t673[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t675 = FSM_fft_64_stage_1_0_t659;
    FSM_fft_64_stage_1_0_t675[FSM_fft_64_stage_1_0_t662 * 32 +: 32] = FSM_fft_64_stage_1_0_t674;
    FSM_fft_64_stage_1_0_t676 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011110;
    FSM_fft_64_stage_1_0_t677 = FSM_fft_64_stage_1_0_t676[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t678 = FSM_fft_64_stage_1_0_t677 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t679 = FSM_fft_64_stage_1_0_t678[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t680 = FSM_fft_64_stage_1_0_t679[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t681 = FSM_fft_64_stage_1_0_t675;
    FSM_fft_64_stage_1_0_t681[FSM_fft_64_stage_1_0_t680 * 32 +: 32] = FSM_fft_64_stage_1_0_t666 - FSM_fft_64_stage_1_0_t672;
    FSM_fft_64_stage_1_0_t682 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011111;
    FSM_fft_64_stage_1_0_t683 = FSM_fft_64_stage_1_0_t682[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t684 = FSM_fft_64_stage_1_0_t683[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t685 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011111;
    FSM_fft_64_stage_1_0_t686 = FSM_fft_64_stage_1_0_t685[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t687 = FSM_fft_64_stage_1_0_t686[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t688 = i_data_in_real[FSM_fft_64_stage_1_0_t687 * 32 +: 32];
    FSM_fft_64_stage_1_0_t689 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011111;
    FSM_fft_64_stage_1_0_t690 = FSM_fft_64_stage_1_0_t689[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t691 = FSM_fft_64_stage_1_0_t690 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t692 = FSM_fft_64_stage_1_0_t691[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t693 = FSM_fft_64_stage_1_0_t692[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t694 = i_data_in_real[FSM_fft_64_stage_1_0_t693 * 32 +: 32];
    FSM_fft_64_stage_1_0_t695 = FSM_fft_64_stage_1_0_t688 + FSM_fft_64_stage_1_0_t694;
    FSM_fft_64_stage_1_0_t696 = FSM_fft_64_stage_1_0_t695[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t697 = FSM_fft_64_stage_1_0_t681;
    FSM_fft_64_stage_1_0_t697[FSM_fft_64_stage_1_0_t684 * 32 +: 32] = FSM_fft_64_stage_1_0_t696;
    FSM_fft_64_stage_1_0_t698 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011111;
    FSM_fft_64_stage_1_0_t699 = FSM_fft_64_stage_1_0_t698[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t700 = FSM_fft_64_stage_1_0_t699 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t701 = FSM_fft_64_stage_1_0_t700[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t702 = FSM_fft_64_stage_1_0_t701[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t703 = FSM_fft_64_stage_1_0_t697;
    FSM_fft_64_stage_1_0_t703[FSM_fft_64_stage_1_0_t702 * 32 +: 32] = FSM_fft_64_stage_1_0_t688 - FSM_fft_64_stage_1_0_t694;
    FSM_fft_64_stage_1_0_t704 = 32'b00000000000000000000000000000010 * 32'b0;
    FSM_fft_64_stage_1_0_t705 = FSM_fft_64_stage_1_0_t704[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t706 = FSM_fft_64_stage_1_0_t705[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t707 = 32'b00000000000000000000000000000010 * 32'b0;
    FSM_fft_64_stage_1_0_t708 = FSM_fft_64_stage_1_0_t707[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t709 = FSM_fft_64_stage_1_0_t708[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t710 = i_data_in_imag[FSM_fft_64_stage_1_0_t709 * 32 +: 32];
    FSM_fft_64_stage_1_0_t711 = 32'b00000000000000000000000000000010 * 32'b0;
    FSM_fft_64_stage_1_0_t712 = FSM_fft_64_stage_1_0_t711[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t713 = FSM_fft_64_stage_1_0_t712 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t714 = FSM_fft_64_stage_1_0_t713[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t715 = FSM_fft_64_stage_1_0_t714[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t716 = i_data_in_imag[FSM_fft_64_stage_1_0_t715 * 32 +: 32];
    FSM_fft_64_stage_1_0_t717 = FSM_fft_64_stage_1_0_t710 + FSM_fft_64_stage_1_0_t716;
    FSM_fft_64_stage_1_0_t718 = FSM_fft_64_stage_1_0_t717[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t719 = 2048'b0;
    FSM_fft_64_stage_1_0_t719[FSM_fft_64_stage_1_0_t706 * 32 +: 32] = FSM_fft_64_stage_1_0_t718;
    FSM_fft_64_stage_1_0_t720 = 32'b00000000000000000000000000000010 * 32'b0;
    FSM_fft_64_stage_1_0_t721 = FSM_fft_64_stage_1_0_t720[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t722 = FSM_fft_64_stage_1_0_t721 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t723 = FSM_fft_64_stage_1_0_t722[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t724 = FSM_fft_64_stage_1_0_t723[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t725 = FSM_fft_64_stage_1_0_t719;
    FSM_fft_64_stage_1_0_t725[FSM_fft_64_stage_1_0_t724 * 32 +: 32] = FSM_fft_64_stage_1_0_t710 - FSM_fft_64_stage_1_0_t716;
    FSM_fft_64_stage_1_0_t726 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t727 = FSM_fft_64_stage_1_0_t726[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t728 = FSM_fft_64_stage_1_0_t727[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t729 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t730 = FSM_fft_64_stage_1_0_t729[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t731 = FSM_fft_64_stage_1_0_t730[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t732 = i_data_in_imag[FSM_fft_64_stage_1_0_t731 * 32 +: 32];
    FSM_fft_64_stage_1_0_t733 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t734 = FSM_fft_64_stage_1_0_t733[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t735 = FSM_fft_64_stage_1_0_t734 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t736 = FSM_fft_64_stage_1_0_t735[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t737 = FSM_fft_64_stage_1_0_t736[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t738 = i_data_in_imag[FSM_fft_64_stage_1_0_t737 * 32 +: 32];
    FSM_fft_64_stage_1_0_t739 = FSM_fft_64_stage_1_0_t732 + FSM_fft_64_stage_1_0_t738;
    FSM_fft_64_stage_1_0_t740 = FSM_fft_64_stage_1_0_t739[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t741 = FSM_fft_64_stage_1_0_t725;
    FSM_fft_64_stage_1_0_t741[FSM_fft_64_stage_1_0_t728 * 32 +: 32] = FSM_fft_64_stage_1_0_t740;
    FSM_fft_64_stage_1_0_t742 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t743 = FSM_fft_64_stage_1_0_t742[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t744 = FSM_fft_64_stage_1_0_t743 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t745 = FSM_fft_64_stage_1_0_t744[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t746 = FSM_fft_64_stage_1_0_t745[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t747 = FSM_fft_64_stage_1_0_t741;
    FSM_fft_64_stage_1_0_t747[FSM_fft_64_stage_1_0_t746 * 32 +: 32] = FSM_fft_64_stage_1_0_t732 - FSM_fft_64_stage_1_0_t738;
    FSM_fft_64_stage_1_0_t748 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_1_0_t749 = FSM_fft_64_stage_1_0_t748[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t750 = FSM_fft_64_stage_1_0_t749[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t751 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_1_0_t752 = FSM_fft_64_stage_1_0_t751[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t753 = FSM_fft_64_stage_1_0_t752[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t754 = i_data_in_imag[FSM_fft_64_stage_1_0_t753 * 32 +: 32];
    FSM_fft_64_stage_1_0_t755 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_1_0_t756 = FSM_fft_64_stage_1_0_t755[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t757 = FSM_fft_64_stage_1_0_t756 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t758 = FSM_fft_64_stage_1_0_t757[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t759 = FSM_fft_64_stage_1_0_t758[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t760 = i_data_in_imag[FSM_fft_64_stage_1_0_t759 * 32 +: 32];
    FSM_fft_64_stage_1_0_t761 = FSM_fft_64_stage_1_0_t754 + FSM_fft_64_stage_1_0_t760;
    FSM_fft_64_stage_1_0_t762 = FSM_fft_64_stage_1_0_t761[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t763 = FSM_fft_64_stage_1_0_t747;
    FSM_fft_64_stage_1_0_t763[FSM_fft_64_stage_1_0_t750 * 32 +: 32] = FSM_fft_64_stage_1_0_t762;
    FSM_fft_64_stage_1_0_t764 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_1_0_t765 = FSM_fft_64_stage_1_0_t764[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t766 = FSM_fft_64_stage_1_0_t765 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t767 = FSM_fft_64_stage_1_0_t766[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t768 = FSM_fft_64_stage_1_0_t767[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t769 = FSM_fft_64_stage_1_0_t763;
    FSM_fft_64_stage_1_0_t769[FSM_fft_64_stage_1_0_t768 * 32 +: 32] = FSM_fft_64_stage_1_0_t754 - FSM_fft_64_stage_1_0_t760;
    FSM_fft_64_stage_1_0_t770 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_1_0_t771 = FSM_fft_64_stage_1_0_t770[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t772 = FSM_fft_64_stage_1_0_t771[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t773 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_1_0_t774 = FSM_fft_64_stage_1_0_t773[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t775 = FSM_fft_64_stage_1_0_t774[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t776 = i_data_in_imag[FSM_fft_64_stage_1_0_t775 * 32 +: 32];
    FSM_fft_64_stage_1_0_t777 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_1_0_t778 = FSM_fft_64_stage_1_0_t777[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t779 = FSM_fft_64_stage_1_0_t778 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t780 = FSM_fft_64_stage_1_0_t779[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t781 = FSM_fft_64_stage_1_0_t780[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t782 = i_data_in_imag[FSM_fft_64_stage_1_0_t781 * 32 +: 32];
    FSM_fft_64_stage_1_0_t783 = FSM_fft_64_stage_1_0_t776 + FSM_fft_64_stage_1_0_t782;
    FSM_fft_64_stage_1_0_t784 = FSM_fft_64_stage_1_0_t783[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t785 = FSM_fft_64_stage_1_0_t769;
    FSM_fft_64_stage_1_0_t785[FSM_fft_64_stage_1_0_t772 * 32 +: 32] = FSM_fft_64_stage_1_0_t784;
    FSM_fft_64_stage_1_0_t786 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_1_0_t787 = FSM_fft_64_stage_1_0_t786[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t788 = FSM_fft_64_stage_1_0_t787 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t789 = FSM_fft_64_stage_1_0_t788[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t790 = FSM_fft_64_stage_1_0_t789[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t791 = FSM_fft_64_stage_1_0_t785;
    FSM_fft_64_stage_1_0_t791[FSM_fft_64_stage_1_0_t790 * 32 +: 32] = FSM_fft_64_stage_1_0_t776 - FSM_fft_64_stage_1_0_t782;
    FSM_fft_64_stage_1_0_t792 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000100;
    FSM_fft_64_stage_1_0_t793 = FSM_fft_64_stage_1_0_t792[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t794 = FSM_fft_64_stage_1_0_t793[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t795 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000100;
    FSM_fft_64_stage_1_0_t796 = FSM_fft_64_stage_1_0_t795[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t797 = FSM_fft_64_stage_1_0_t796[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t798 = i_data_in_imag[FSM_fft_64_stage_1_0_t797 * 32 +: 32];
    FSM_fft_64_stage_1_0_t799 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000100;
    FSM_fft_64_stage_1_0_t800 = FSM_fft_64_stage_1_0_t799[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t801 = FSM_fft_64_stage_1_0_t800 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t802 = FSM_fft_64_stage_1_0_t801[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t803 = FSM_fft_64_stage_1_0_t802[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t804 = i_data_in_imag[FSM_fft_64_stage_1_0_t803 * 32 +: 32];
    FSM_fft_64_stage_1_0_t805 = FSM_fft_64_stage_1_0_t798 + FSM_fft_64_stage_1_0_t804;
    FSM_fft_64_stage_1_0_t806 = FSM_fft_64_stage_1_0_t805[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t807 = FSM_fft_64_stage_1_0_t791;
    FSM_fft_64_stage_1_0_t807[FSM_fft_64_stage_1_0_t794 * 32 +: 32] = FSM_fft_64_stage_1_0_t806;
    FSM_fft_64_stage_1_0_t808 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000100;
    FSM_fft_64_stage_1_0_t809 = FSM_fft_64_stage_1_0_t808[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t810 = FSM_fft_64_stage_1_0_t809 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t811 = FSM_fft_64_stage_1_0_t810[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t812 = FSM_fft_64_stage_1_0_t811[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t813 = FSM_fft_64_stage_1_0_t807;
    FSM_fft_64_stage_1_0_t813[FSM_fft_64_stage_1_0_t812 * 32 +: 32] = FSM_fft_64_stage_1_0_t798 - FSM_fft_64_stage_1_0_t804;
    FSM_fft_64_stage_1_0_t814 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000101;
    FSM_fft_64_stage_1_0_t815 = FSM_fft_64_stage_1_0_t814[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t816 = FSM_fft_64_stage_1_0_t815[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t817 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000101;
    FSM_fft_64_stage_1_0_t818 = FSM_fft_64_stage_1_0_t817[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t819 = FSM_fft_64_stage_1_0_t818[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t820 = i_data_in_imag[FSM_fft_64_stage_1_0_t819 * 32 +: 32];
    FSM_fft_64_stage_1_0_t821 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000101;
    FSM_fft_64_stage_1_0_t822 = FSM_fft_64_stage_1_0_t821[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t823 = FSM_fft_64_stage_1_0_t822 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t824 = FSM_fft_64_stage_1_0_t823[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t825 = FSM_fft_64_stage_1_0_t824[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t826 = i_data_in_imag[FSM_fft_64_stage_1_0_t825 * 32 +: 32];
    FSM_fft_64_stage_1_0_t827 = FSM_fft_64_stage_1_0_t820 + FSM_fft_64_stage_1_0_t826;
    FSM_fft_64_stage_1_0_t828 = FSM_fft_64_stage_1_0_t827[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t829 = FSM_fft_64_stage_1_0_t813;
    FSM_fft_64_stage_1_0_t829[FSM_fft_64_stage_1_0_t816 * 32 +: 32] = FSM_fft_64_stage_1_0_t828;
    FSM_fft_64_stage_1_0_t830 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000101;
    FSM_fft_64_stage_1_0_t831 = FSM_fft_64_stage_1_0_t830[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t832 = FSM_fft_64_stage_1_0_t831 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t833 = FSM_fft_64_stage_1_0_t832[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t834 = FSM_fft_64_stage_1_0_t833[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t835 = FSM_fft_64_stage_1_0_t829;
    FSM_fft_64_stage_1_0_t835[FSM_fft_64_stage_1_0_t834 * 32 +: 32] = FSM_fft_64_stage_1_0_t820 - FSM_fft_64_stage_1_0_t826;
    FSM_fft_64_stage_1_0_t836 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000110;
    FSM_fft_64_stage_1_0_t837 = FSM_fft_64_stage_1_0_t836[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t838 = FSM_fft_64_stage_1_0_t837[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t839 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000110;
    FSM_fft_64_stage_1_0_t840 = FSM_fft_64_stage_1_0_t839[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t841 = FSM_fft_64_stage_1_0_t840[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t842 = i_data_in_imag[FSM_fft_64_stage_1_0_t841 * 32 +: 32];
    FSM_fft_64_stage_1_0_t843 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000110;
    FSM_fft_64_stage_1_0_t844 = FSM_fft_64_stage_1_0_t843[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t845 = FSM_fft_64_stage_1_0_t844 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t846 = FSM_fft_64_stage_1_0_t845[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t847 = FSM_fft_64_stage_1_0_t846[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t848 = i_data_in_imag[FSM_fft_64_stage_1_0_t847 * 32 +: 32];
    FSM_fft_64_stage_1_0_t849 = FSM_fft_64_stage_1_0_t842 + FSM_fft_64_stage_1_0_t848;
    FSM_fft_64_stage_1_0_t850 = FSM_fft_64_stage_1_0_t849[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t851 = FSM_fft_64_stage_1_0_t835;
    FSM_fft_64_stage_1_0_t851[FSM_fft_64_stage_1_0_t838 * 32 +: 32] = FSM_fft_64_stage_1_0_t850;
    FSM_fft_64_stage_1_0_t852 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000110;
    FSM_fft_64_stage_1_0_t853 = FSM_fft_64_stage_1_0_t852[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t854 = FSM_fft_64_stage_1_0_t853 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t855 = FSM_fft_64_stage_1_0_t854[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t856 = FSM_fft_64_stage_1_0_t855[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t857 = FSM_fft_64_stage_1_0_t851;
    FSM_fft_64_stage_1_0_t857[FSM_fft_64_stage_1_0_t856 * 32 +: 32] = FSM_fft_64_stage_1_0_t842 - FSM_fft_64_stage_1_0_t848;
    FSM_fft_64_stage_1_0_t858 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000111;
    FSM_fft_64_stage_1_0_t859 = FSM_fft_64_stage_1_0_t858[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t860 = FSM_fft_64_stage_1_0_t859[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t861 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000111;
    FSM_fft_64_stage_1_0_t862 = FSM_fft_64_stage_1_0_t861[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t863 = FSM_fft_64_stage_1_0_t862[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t864 = i_data_in_imag[FSM_fft_64_stage_1_0_t863 * 32 +: 32];
    FSM_fft_64_stage_1_0_t865 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000111;
    FSM_fft_64_stage_1_0_t866 = FSM_fft_64_stage_1_0_t865[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t867 = FSM_fft_64_stage_1_0_t866 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t868 = FSM_fft_64_stage_1_0_t867[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t869 = FSM_fft_64_stage_1_0_t868[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t870 = i_data_in_imag[FSM_fft_64_stage_1_0_t869 * 32 +: 32];
    FSM_fft_64_stage_1_0_t871 = FSM_fft_64_stage_1_0_t864 + FSM_fft_64_stage_1_0_t870;
    FSM_fft_64_stage_1_0_t872 = FSM_fft_64_stage_1_0_t871[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t873 = FSM_fft_64_stage_1_0_t857;
    FSM_fft_64_stage_1_0_t873[FSM_fft_64_stage_1_0_t860 * 32 +: 32] = FSM_fft_64_stage_1_0_t872;
    FSM_fft_64_stage_1_0_t874 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000000111;
    FSM_fft_64_stage_1_0_t875 = FSM_fft_64_stage_1_0_t874[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t876 = FSM_fft_64_stage_1_0_t875 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t877 = FSM_fft_64_stage_1_0_t876[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t878 = FSM_fft_64_stage_1_0_t877[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t879 = FSM_fft_64_stage_1_0_t873;
    FSM_fft_64_stage_1_0_t879[FSM_fft_64_stage_1_0_t878 * 32 +: 32] = FSM_fft_64_stage_1_0_t864 - FSM_fft_64_stage_1_0_t870;
    FSM_fft_64_stage_1_0_t880 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001000;
    FSM_fft_64_stage_1_0_t881 = FSM_fft_64_stage_1_0_t880[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t882 = FSM_fft_64_stage_1_0_t881[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t883 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001000;
    FSM_fft_64_stage_1_0_t884 = FSM_fft_64_stage_1_0_t883[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t885 = FSM_fft_64_stage_1_0_t884[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t886 = i_data_in_imag[FSM_fft_64_stage_1_0_t885 * 32 +: 32];
    FSM_fft_64_stage_1_0_t887 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001000;
    FSM_fft_64_stage_1_0_t888 = FSM_fft_64_stage_1_0_t887[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t889 = FSM_fft_64_stage_1_0_t888 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t890 = FSM_fft_64_stage_1_0_t889[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t891 = FSM_fft_64_stage_1_0_t890[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t892 = i_data_in_imag[FSM_fft_64_stage_1_0_t891 * 32 +: 32];
    FSM_fft_64_stage_1_0_t893 = FSM_fft_64_stage_1_0_t886 + FSM_fft_64_stage_1_0_t892;
    FSM_fft_64_stage_1_0_t894 = FSM_fft_64_stage_1_0_t893[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t895 = FSM_fft_64_stage_1_0_t879;
    FSM_fft_64_stage_1_0_t895[FSM_fft_64_stage_1_0_t882 * 32 +: 32] = FSM_fft_64_stage_1_0_t894;
    FSM_fft_64_stage_1_0_t896 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001000;
    FSM_fft_64_stage_1_0_t897 = FSM_fft_64_stage_1_0_t896[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t898 = FSM_fft_64_stage_1_0_t897 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t899 = FSM_fft_64_stage_1_0_t898[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t900 = FSM_fft_64_stage_1_0_t899[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t901 = FSM_fft_64_stage_1_0_t895;
    FSM_fft_64_stage_1_0_t901[FSM_fft_64_stage_1_0_t900 * 32 +: 32] = FSM_fft_64_stage_1_0_t886 - FSM_fft_64_stage_1_0_t892;
    FSM_fft_64_stage_1_0_t902 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001001;
    FSM_fft_64_stage_1_0_t903 = FSM_fft_64_stage_1_0_t902[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t904 = FSM_fft_64_stage_1_0_t903[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t905 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001001;
    FSM_fft_64_stage_1_0_t906 = FSM_fft_64_stage_1_0_t905[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t907 = FSM_fft_64_stage_1_0_t906[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t908 = i_data_in_imag[FSM_fft_64_stage_1_0_t907 * 32 +: 32];
    FSM_fft_64_stage_1_0_t909 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001001;
    FSM_fft_64_stage_1_0_t910 = FSM_fft_64_stage_1_0_t909[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t911 = FSM_fft_64_stage_1_0_t910 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t912 = FSM_fft_64_stage_1_0_t911[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t913 = FSM_fft_64_stage_1_0_t912[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t914 = i_data_in_imag[FSM_fft_64_stage_1_0_t913 * 32 +: 32];
    FSM_fft_64_stage_1_0_t915 = FSM_fft_64_stage_1_0_t908 + FSM_fft_64_stage_1_0_t914;
    FSM_fft_64_stage_1_0_t916 = FSM_fft_64_stage_1_0_t915[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t917 = FSM_fft_64_stage_1_0_t901;
    FSM_fft_64_stage_1_0_t917[FSM_fft_64_stage_1_0_t904 * 32 +: 32] = FSM_fft_64_stage_1_0_t916;
    FSM_fft_64_stage_1_0_t918 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001001;
    FSM_fft_64_stage_1_0_t919 = FSM_fft_64_stage_1_0_t918[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t920 = FSM_fft_64_stage_1_0_t919 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t921 = FSM_fft_64_stage_1_0_t920[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t922 = FSM_fft_64_stage_1_0_t921[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t923 = FSM_fft_64_stage_1_0_t917;
    FSM_fft_64_stage_1_0_t923[FSM_fft_64_stage_1_0_t922 * 32 +: 32] = FSM_fft_64_stage_1_0_t908 - FSM_fft_64_stage_1_0_t914;
    FSM_fft_64_stage_1_0_t924 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001010;
    FSM_fft_64_stage_1_0_t925 = FSM_fft_64_stage_1_0_t924[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t926 = FSM_fft_64_stage_1_0_t925[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t927 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001010;
    FSM_fft_64_stage_1_0_t928 = FSM_fft_64_stage_1_0_t927[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t929 = FSM_fft_64_stage_1_0_t928[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t930 = i_data_in_imag[FSM_fft_64_stage_1_0_t929 * 32 +: 32];
    FSM_fft_64_stage_1_0_t931 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001010;
    FSM_fft_64_stage_1_0_t932 = FSM_fft_64_stage_1_0_t931[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t933 = FSM_fft_64_stage_1_0_t932 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t934 = FSM_fft_64_stage_1_0_t933[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t935 = FSM_fft_64_stage_1_0_t934[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t936 = i_data_in_imag[FSM_fft_64_stage_1_0_t935 * 32 +: 32];
    FSM_fft_64_stage_1_0_t937 = FSM_fft_64_stage_1_0_t930 + FSM_fft_64_stage_1_0_t936;
    FSM_fft_64_stage_1_0_t938 = FSM_fft_64_stage_1_0_t937[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t939 = FSM_fft_64_stage_1_0_t923;
    FSM_fft_64_stage_1_0_t939[FSM_fft_64_stage_1_0_t926 * 32 +: 32] = FSM_fft_64_stage_1_0_t938;
    FSM_fft_64_stage_1_0_t940 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001010;
    FSM_fft_64_stage_1_0_t941 = FSM_fft_64_stage_1_0_t940[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t942 = FSM_fft_64_stage_1_0_t941 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t943 = FSM_fft_64_stage_1_0_t942[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t944 = FSM_fft_64_stage_1_0_t943[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t945 = FSM_fft_64_stage_1_0_t939;
    FSM_fft_64_stage_1_0_t945[FSM_fft_64_stage_1_0_t944 * 32 +: 32] = FSM_fft_64_stage_1_0_t930 - FSM_fft_64_stage_1_0_t936;
    FSM_fft_64_stage_1_0_t946 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001011;
    FSM_fft_64_stage_1_0_t947 = FSM_fft_64_stage_1_0_t946[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t948 = FSM_fft_64_stage_1_0_t947[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t949 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001011;
    FSM_fft_64_stage_1_0_t950 = FSM_fft_64_stage_1_0_t949[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t951 = FSM_fft_64_stage_1_0_t950[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t952 = i_data_in_imag[FSM_fft_64_stage_1_0_t951 * 32 +: 32];
    FSM_fft_64_stage_1_0_t953 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001011;
    FSM_fft_64_stage_1_0_t954 = FSM_fft_64_stage_1_0_t953[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t955 = FSM_fft_64_stage_1_0_t954 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t956 = FSM_fft_64_stage_1_0_t955[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t957 = FSM_fft_64_stage_1_0_t956[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t958 = i_data_in_imag[FSM_fft_64_stage_1_0_t957 * 32 +: 32];
    FSM_fft_64_stage_1_0_t959 = FSM_fft_64_stage_1_0_t952 + FSM_fft_64_stage_1_0_t958;
    FSM_fft_64_stage_1_0_t960 = FSM_fft_64_stage_1_0_t959[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t961 = FSM_fft_64_stage_1_0_t945;
    FSM_fft_64_stage_1_0_t961[FSM_fft_64_stage_1_0_t948 * 32 +: 32] = FSM_fft_64_stage_1_0_t960;
    FSM_fft_64_stage_1_0_t962 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001011;
    FSM_fft_64_stage_1_0_t963 = FSM_fft_64_stage_1_0_t962[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t964 = FSM_fft_64_stage_1_0_t963 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t965 = FSM_fft_64_stage_1_0_t964[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t966 = FSM_fft_64_stage_1_0_t965[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t967 = FSM_fft_64_stage_1_0_t961;
    FSM_fft_64_stage_1_0_t967[FSM_fft_64_stage_1_0_t966 * 32 +: 32] = FSM_fft_64_stage_1_0_t952 - FSM_fft_64_stage_1_0_t958;
    FSM_fft_64_stage_1_0_t968 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001100;
    FSM_fft_64_stage_1_0_t969 = FSM_fft_64_stage_1_0_t968[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t970 = FSM_fft_64_stage_1_0_t969[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t971 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001100;
    FSM_fft_64_stage_1_0_t972 = FSM_fft_64_stage_1_0_t971[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t973 = FSM_fft_64_stage_1_0_t972[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t974 = i_data_in_imag[FSM_fft_64_stage_1_0_t973 * 32 +: 32];
    FSM_fft_64_stage_1_0_t975 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001100;
    FSM_fft_64_stage_1_0_t976 = FSM_fft_64_stage_1_0_t975[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t977 = FSM_fft_64_stage_1_0_t976 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t978 = FSM_fft_64_stage_1_0_t977[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t979 = FSM_fft_64_stage_1_0_t978[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t980 = i_data_in_imag[FSM_fft_64_stage_1_0_t979 * 32 +: 32];
    FSM_fft_64_stage_1_0_t981 = FSM_fft_64_stage_1_0_t974 + FSM_fft_64_stage_1_0_t980;
    FSM_fft_64_stage_1_0_t982 = FSM_fft_64_stage_1_0_t981[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t983 = FSM_fft_64_stage_1_0_t967;
    FSM_fft_64_stage_1_0_t983[FSM_fft_64_stage_1_0_t970 * 32 +: 32] = FSM_fft_64_stage_1_0_t982;
    FSM_fft_64_stage_1_0_t984 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001100;
    FSM_fft_64_stage_1_0_t985 = FSM_fft_64_stage_1_0_t984[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t986 = FSM_fft_64_stage_1_0_t985 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t987 = FSM_fft_64_stage_1_0_t986[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t988 = FSM_fft_64_stage_1_0_t987[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t989 = FSM_fft_64_stage_1_0_t983;
    FSM_fft_64_stage_1_0_t989[FSM_fft_64_stage_1_0_t988 * 32 +: 32] = FSM_fft_64_stage_1_0_t974 - FSM_fft_64_stage_1_0_t980;
    FSM_fft_64_stage_1_0_t990 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001101;
    FSM_fft_64_stage_1_0_t991 = FSM_fft_64_stage_1_0_t990[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t992 = FSM_fft_64_stage_1_0_t991[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t993 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001101;
    FSM_fft_64_stage_1_0_t994 = FSM_fft_64_stage_1_0_t993[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t995 = FSM_fft_64_stage_1_0_t994[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t996 = i_data_in_imag[FSM_fft_64_stage_1_0_t995 * 32 +: 32];
    FSM_fft_64_stage_1_0_t997 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001101;
    FSM_fft_64_stage_1_0_t998 = FSM_fft_64_stage_1_0_t997[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t999 = FSM_fft_64_stage_1_0_t998 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1000 = FSM_fft_64_stage_1_0_t999[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1001 = FSM_fft_64_stage_1_0_t1000[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1002 = i_data_in_imag[FSM_fft_64_stage_1_0_t1001 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1003 = FSM_fft_64_stage_1_0_t996 + FSM_fft_64_stage_1_0_t1002;
    FSM_fft_64_stage_1_0_t1004 = FSM_fft_64_stage_1_0_t1003[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1005 = FSM_fft_64_stage_1_0_t989;
    FSM_fft_64_stage_1_0_t1005[FSM_fft_64_stage_1_0_t992 * 32 +: 32] = FSM_fft_64_stage_1_0_t1004;
    FSM_fft_64_stage_1_0_t1006 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001101;
    FSM_fft_64_stage_1_0_t1007 = FSM_fft_64_stage_1_0_t1006[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1008 = FSM_fft_64_stage_1_0_t1007 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1009 = FSM_fft_64_stage_1_0_t1008[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1010 = FSM_fft_64_stage_1_0_t1009[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1011 = FSM_fft_64_stage_1_0_t1005;
    FSM_fft_64_stage_1_0_t1011[FSM_fft_64_stage_1_0_t1010 * 32 +: 32] = FSM_fft_64_stage_1_0_t996 - FSM_fft_64_stage_1_0_t1002;
    FSM_fft_64_stage_1_0_t1012 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001110;
    FSM_fft_64_stage_1_0_t1013 = FSM_fft_64_stage_1_0_t1012[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1014 = FSM_fft_64_stage_1_0_t1013[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1015 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001110;
    FSM_fft_64_stage_1_0_t1016 = FSM_fft_64_stage_1_0_t1015[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1017 = FSM_fft_64_stage_1_0_t1016[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1018 = i_data_in_imag[FSM_fft_64_stage_1_0_t1017 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1019 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001110;
    FSM_fft_64_stage_1_0_t1020 = FSM_fft_64_stage_1_0_t1019[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1021 = FSM_fft_64_stage_1_0_t1020 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1022 = FSM_fft_64_stage_1_0_t1021[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1023 = FSM_fft_64_stage_1_0_t1022[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1024 = i_data_in_imag[FSM_fft_64_stage_1_0_t1023 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1025 = FSM_fft_64_stage_1_0_t1018 + FSM_fft_64_stage_1_0_t1024;
    FSM_fft_64_stage_1_0_t1026 = FSM_fft_64_stage_1_0_t1025[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1027 = FSM_fft_64_stage_1_0_t1011;
    FSM_fft_64_stage_1_0_t1027[FSM_fft_64_stage_1_0_t1014 * 32 +: 32] = FSM_fft_64_stage_1_0_t1026;
    FSM_fft_64_stage_1_0_t1028 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001110;
    FSM_fft_64_stage_1_0_t1029 = FSM_fft_64_stage_1_0_t1028[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1030 = FSM_fft_64_stage_1_0_t1029 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1031 = FSM_fft_64_stage_1_0_t1030[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1032 = FSM_fft_64_stage_1_0_t1031[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1033 = FSM_fft_64_stage_1_0_t1027;
    FSM_fft_64_stage_1_0_t1033[FSM_fft_64_stage_1_0_t1032 * 32 +: 32] = FSM_fft_64_stage_1_0_t1018 - FSM_fft_64_stage_1_0_t1024;
    FSM_fft_64_stage_1_0_t1034 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001111;
    FSM_fft_64_stage_1_0_t1035 = FSM_fft_64_stage_1_0_t1034[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1036 = FSM_fft_64_stage_1_0_t1035[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1037 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001111;
    FSM_fft_64_stage_1_0_t1038 = FSM_fft_64_stage_1_0_t1037[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1039 = FSM_fft_64_stage_1_0_t1038[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1040 = i_data_in_imag[FSM_fft_64_stage_1_0_t1039 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1041 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001111;
    FSM_fft_64_stage_1_0_t1042 = FSM_fft_64_stage_1_0_t1041[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1043 = FSM_fft_64_stage_1_0_t1042 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1044 = FSM_fft_64_stage_1_0_t1043[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1045 = FSM_fft_64_stage_1_0_t1044[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1046 = i_data_in_imag[FSM_fft_64_stage_1_0_t1045 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1047 = FSM_fft_64_stage_1_0_t1040 + FSM_fft_64_stage_1_0_t1046;
    FSM_fft_64_stage_1_0_t1048 = FSM_fft_64_stage_1_0_t1047[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1049 = FSM_fft_64_stage_1_0_t1033;
    FSM_fft_64_stage_1_0_t1049[FSM_fft_64_stage_1_0_t1036 * 32 +: 32] = FSM_fft_64_stage_1_0_t1048;
    FSM_fft_64_stage_1_0_t1050 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000001111;
    FSM_fft_64_stage_1_0_t1051 = FSM_fft_64_stage_1_0_t1050[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1052 = FSM_fft_64_stage_1_0_t1051 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1053 = FSM_fft_64_stage_1_0_t1052[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1054 = FSM_fft_64_stage_1_0_t1053[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1055 = FSM_fft_64_stage_1_0_t1049;
    FSM_fft_64_stage_1_0_t1055[FSM_fft_64_stage_1_0_t1054 * 32 +: 32] = FSM_fft_64_stage_1_0_t1040 - FSM_fft_64_stage_1_0_t1046;
    FSM_fft_64_stage_1_0_t1056 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010000;
    FSM_fft_64_stage_1_0_t1057 = FSM_fft_64_stage_1_0_t1056[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1058 = FSM_fft_64_stage_1_0_t1057[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1059 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010000;
    FSM_fft_64_stage_1_0_t1060 = FSM_fft_64_stage_1_0_t1059[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1061 = FSM_fft_64_stage_1_0_t1060[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1062 = i_data_in_imag[FSM_fft_64_stage_1_0_t1061 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1063 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010000;
    FSM_fft_64_stage_1_0_t1064 = FSM_fft_64_stage_1_0_t1063[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1065 = FSM_fft_64_stage_1_0_t1064 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1066 = FSM_fft_64_stage_1_0_t1065[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1067 = FSM_fft_64_stage_1_0_t1066[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1068 = i_data_in_imag[FSM_fft_64_stage_1_0_t1067 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1069 = FSM_fft_64_stage_1_0_t1062 + FSM_fft_64_stage_1_0_t1068;
    FSM_fft_64_stage_1_0_t1070 = FSM_fft_64_stage_1_0_t1069[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1071 = FSM_fft_64_stage_1_0_t1055;
    FSM_fft_64_stage_1_0_t1071[FSM_fft_64_stage_1_0_t1058 * 32 +: 32] = FSM_fft_64_stage_1_0_t1070;
    FSM_fft_64_stage_1_0_t1072 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010000;
    FSM_fft_64_stage_1_0_t1073 = FSM_fft_64_stage_1_0_t1072[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1074 = FSM_fft_64_stage_1_0_t1073 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1075 = FSM_fft_64_stage_1_0_t1074[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1076 = FSM_fft_64_stage_1_0_t1075[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1077 = FSM_fft_64_stage_1_0_t1071;
    FSM_fft_64_stage_1_0_t1077[FSM_fft_64_stage_1_0_t1076 * 32 +: 32] = FSM_fft_64_stage_1_0_t1062 - FSM_fft_64_stage_1_0_t1068;
    FSM_fft_64_stage_1_0_t1078 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010001;
    FSM_fft_64_stage_1_0_t1079 = FSM_fft_64_stage_1_0_t1078[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1080 = FSM_fft_64_stage_1_0_t1079[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1081 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010001;
    FSM_fft_64_stage_1_0_t1082 = FSM_fft_64_stage_1_0_t1081[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1083 = FSM_fft_64_stage_1_0_t1082[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1084 = i_data_in_imag[FSM_fft_64_stage_1_0_t1083 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1085 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010001;
    FSM_fft_64_stage_1_0_t1086 = FSM_fft_64_stage_1_0_t1085[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1087 = FSM_fft_64_stage_1_0_t1086 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1088 = FSM_fft_64_stage_1_0_t1087[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1089 = FSM_fft_64_stage_1_0_t1088[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1090 = i_data_in_imag[FSM_fft_64_stage_1_0_t1089 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1091 = FSM_fft_64_stage_1_0_t1084 + FSM_fft_64_stage_1_0_t1090;
    FSM_fft_64_stage_1_0_t1092 = FSM_fft_64_stage_1_0_t1091[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1093 = FSM_fft_64_stage_1_0_t1077;
    FSM_fft_64_stage_1_0_t1093[FSM_fft_64_stage_1_0_t1080 * 32 +: 32] = FSM_fft_64_stage_1_0_t1092;
    FSM_fft_64_stage_1_0_t1094 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010001;
    FSM_fft_64_stage_1_0_t1095 = FSM_fft_64_stage_1_0_t1094[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1096 = FSM_fft_64_stage_1_0_t1095 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1097 = FSM_fft_64_stage_1_0_t1096[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1098 = FSM_fft_64_stage_1_0_t1097[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1099 = FSM_fft_64_stage_1_0_t1093;
    FSM_fft_64_stage_1_0_t1099[FSM_fft_64_stage_1_0_t1098 * 32 +: 32] = FSM_fft_64_stage_1_0_t1084 - FSM_fft_64_stage_1_0_t1090;
    FSM_fft_64_stage_1_0_t1100 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010010;
    FSM_fft_64_stage_1_0_t1101 = FSM_fft_64_stage_1_0_t1100[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1102 = FSM_fft_64_stage_1_0_t1101[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1103 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010010;
    FSM_fft_64_stage_1_0_t1104 = FSM_fft_64_stage_1_0_t1103[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1105 = FSM_fft_64_stage_1_0_t1104[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1106 = i_data_in_imag[FSM_fft_64_stage_1_0_t1105 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1107 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010010;
    FSM_fft_64_stage_1_0_t1108 = FSM_fft_64_stage_1_0_t1107[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1109 = FSM_fft_64_stage_1_0_t1108 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1110 = FSM_fft_64_stage_1_0_t1109[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1111 = FSM_fft_64_stage_1_0_t1110[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1112 = i_data_in_imag[FSM_fft_64_stage_1_0_t1111 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1113 = FSM_fft_64_stage_1_0_t1106 + FSM_fft_64_stage_1_0_t1112;
    FSM_fft_64_stage_1_0_t1114 = FSM_fft_64_stage_1_0_t1113[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1115 = FSM_fft_64_stage_1_0_t1099;
    FSM_fft_64_stage_1_0_t1115[FSM_fft_64_stage_1_0_t1102 * 32 +: 32] = FSM_fft_64_stage_1_0_t1114;
    FSM_fft_64_stage_1_0_t1116 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010010;
    FSM_fft_64_stage_1_0_t1117 = FSM_fft_64_stage_1_0_t1116[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1118 = FSM_fft_64_stage_1_0_t1117 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1119 = FSM_fft_64_stage_1_0_t1118[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1120 = FSM_fft_64_stage_1_0_t1119[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1121 = FSM_fft_64_stage_1_0_t1115;
    FSM_fft_64_stage_1_0_t1121[FSM_fft_64_stage_1_0_t1120 * 32 +: 32] = FSM_fft_64_stage_1_0_t1106 - FSM_fft_64_stage_1_0_t1112;
    FSM_fft_64_stage_1_0_t1122 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010011;
    FSM_fft_64_stage_1_0_t1123 = FSM_fft_64_stage_1_0_t1122[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1124 = FSM_fft_64_stage_1_0_t1123[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1125 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010011;
    FSM_fft_64_stage_1_0_t1126 = FSM_fft_64_stage_1_0_t1125[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1127 = FSM_fft_64_stage_1_0_t1126[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1128 = i_data_in_imag[FSM_fft_64_stage_1_0_t1127 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1129 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010011;
    FSM_fft_64_stage_1_0_t1130 = FSM_fft_64_stage_1_0_t1129[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1131 = FSM_fft_64_stage_1_0_t1130 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1132 = FSM_fft_64_stage_1_0_t1131[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1133 = FSM_fft_64_stage_1_0_t1132[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1134 = i_data_in_imag[FSM_fft_64_stage_1_0_t1133 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1135 = FSM_fft_64_stage_1_0_t1128 + FSM_fft_64_stage_1_0_t1134;
    FSM_fft_64_stage_1_0_t1136 = FSM_fft_64_stage_1_0_t1135[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1137 = FSM_fft_64_stage_1_0_t1121;
    FSM_fft_64_stage_1_0_t1137[FSM_fft_64_stage_1_0_t1124 * 32 +: 32] = FSM_fft_64_stage_1_0_t1136;
    FSM_fft_64_stage_1_0_t1138 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010011;
    FSM_fft_64_stage_1_0_t1139 = FSM_fft_64_stage_1_0_t1138[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1140 = FSM_fft_64_stage_1_0_t1139 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1141 = FSM_fft_64_stage_1_0_t1140[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1142 = FSM_fft_64_stage_1_0_t1141[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1143 = FSM_fft_64_stage_1_0_t1137;
    FSM_fft_64_stage_1_0_t1143[FSM_fft_64_stage_1_0_t1142 * 32 +: 32] = FSM_fft_64_stage_1_0_t1128 - FSM_fft_64_stage_1_0_t1134;
    FSM_fft_64_stage_1_0_t1144 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010100;
    FSM_fft_64_stage_1_0_t1145 = FSM_fft_64_stage_1_0_t1144[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1146 = FSM_fft_64_stage_1_0_t1145[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1147 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010100;
    FSM_fft_64_stage_1_0_t1148 = FSM_fft_64_stage_1_0_t1147[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1149 = FSM_fft_64_stage_1_0_t1148[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1150 = i_data_in_imag[FSM_fft_64_stage_1_0_t1149 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1151 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010100;
    FSM_fft_64_stage_1_0_t1152 = FSM_fft_64_stage_1_0_t1151[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1153 = FSM_fft_64_stage_1_0_t1152 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1154 = FSM_fft_64_stage_1_0_t1153[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1155 = FSM_fft_64_stage_1_0_t1154[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1156 = i_data_in_imag[FSM_fft_64_stage_1_0_t1155 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1157 = FSM_fft_64_stage_1_0_t1150 + FSM_fft_64_stage_1_0_t1156;
    FSM_fft_64_stage_1_0_t1158 = FSM_fft_64_stage_1_0_t1157[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1159 = FSM_fft_64_stage_1_0_t1143;
    FSM_fft_64_stage_1_0_t1159[FSM_fft_64_stage_1_0_t1146 * 32 +: 32] = FSM_fft_64_stage_1_0_t1158;
    FSM_fft_64_stage_1_0_t1160 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010100;
    FSM_fft_64_stage_1_0_t1161 = FSM_fft_64_stage_1_0_t1160[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1162 = FSM_fft_64_stage_1_0_t1161 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1163 = FSM_fft_64_stage_1_0_t1162[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1164 = FSM_fft_64_stage_1_0_t1163[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1165 = FSM_fft_64_stage_1_0_t1159;
    FSM_fft_64_stage_1_0_t1165[FSM_fft_64_stage_1_0_t1164 * 32 +: 32] = FSM_fft_64_stage_1_0_t1150 - FSM_fft_64_stage_1_0_t1156;
    FSM_fft_64_stage_1_0_t1166 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010101;
    FSM_fft_64_stage_1_0_t1167 = FSM_fft_64_stage_1_0_t1166[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1168 = FSM_fft_64_stage_1_0_t1167[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1169 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010101;
    FSM_fft_64_stage_1_0_t1170 = FSM_fft_64_stage_1_0_t1169[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1171 = FSM_fft_64_stage_1_0_t1170[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1172 = i_data_in_imag[FSM_fft_64_stage_1_0_t1171 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1173 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010101;
    FSM_fft_64_stage_1_0_t1174 = FSM_fft_64_stage_1_0_t1173[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1175 = FSM_fft_64_stage_1_0_t1174 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1176 = FSM_fft_64_stage_1_0_t1175[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1177 = FSM_fft_64_stage_1_0_t1176[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1178 = i_data_in_imag[FSM_fft_64_stage_1_0_t1177 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1179 = FSM_fft_64_stage_1_0_t1172 + FSM_fft_64_stage_1_0_t1178;
    FSM_fft_64_stage_1_0_t1180 = FSM_fft_64_stage_1_0_t1179[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1181 = FSM_fft_64_stage_1_0_t1165;
    FSM_fft_64_stage_1_0_t1181[FSM_fft_64_stage_1_0_t1168 * 32 +: 32] = FSM_fft_64_stage_1_0_t1180;
    FSM_fft_64_stage_1_0_t1182 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010101;
    FSM_fft_64_stage_1_0_t1183 = FSM_fft_64_stage_1_0_t1182[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1184 = FSM_fft_64_stage_1_0_t1183 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1185 = FSM_fft_64_stage_1_0_t1184[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1186 = FSM_fft_64_stage_1_0_t1185[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1187 = FSM_fft_64_stage_1_0_t1181;
    FSM_fft_64_stage_1_0_t1187[FSM_fft_64_stage_1_0_t1186 * 32 +: 32] = FSM_fft_64_stage_1_0_t1172 - FSM_fft_64_stage_1_0_t1178;
    FSM_fft_64_stage_1_0_t1188 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010110;
    FSM_fft_64_stage_1_0_t1189 = FSM_fft_64_stage_1_0_t1188[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1190 = FSM_fft_64_stage_1_0_t1189[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1191 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010110;
    FSM_fft_64_stage_1_0_t1192 = FSM_fft_64_stage_1_0_t1191[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1193 = FSM_fft_64_stage_1_0_t1192[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1194 = i_data_in_imag[FSM_fft_64_stage_1_0_t1193 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1195 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010110;
    FSM_fft_64_stage_1_0_t1196 = FSM_fft_64_stage_1_0_t1195[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1197 = FSM_fft_64_stage_1_0_t1196 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1198 = FSM_fft_64_stage_1_0_t1197[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1199 = FSM_fft_64_stage_1_0_t1198[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1200 = i_data_in_imag[FSM_fft_64_stage_1_0_t1199 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1201 = FSM_fft_64_stage_1_0_t1194 + FSM_fft_64_stage_1_0_t1200;
    FSM_fft_64_stage_1_0_t1202 = FSM_fft_64_stage_1_0_t1201[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1203 = FSM_fft_64_stage_1_0_t1187;
    FSM_fft_64_stage_1_0_t1203[FSM_fft_64_stage_1_0_t1190 * 32 +: 32] = FSM_fft_64_stage_1_0_t1202;
    FSM_fft_64_stage_1_0_t1204 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010110;
    FSM_fft_64_stage_1_0_t1205 = FSM_fft_64_stage_1_0_t1204[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1206 = FSM_fft_64_stage_1_0_t1205 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1207 = FSM_fft_64_stage_1_0_t1206[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1208 = FSM_fft_64_stage_1_0_t1207[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1209 = FSM_fft_64_stage_1_0_t1203;
    FSM_fft_64_stage_1_0_t1209[FSM_fft_64_stage_1_0_t1208 * 32 +: 32] = FSM_fft_64_stage_1_0_t1194 - FSM_fft_64_stage_1_0_t1200;
    FSM_fft_64_stage_1_0_t1210 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010111;
    FSM_fft_64_stage_1_0_t1211 = FSM_fft_64_stage_1_0_t1210[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1212 = FSM_fft_64_stage_1_0_t1211[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1213 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010111;
    FSM_fft_64_stage_1_0_t1214 = FSM_fft_64_stage_1_0_t1213[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1215 = FSM_fft_64_stage_1_0_t1214[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1216 = i_data_in_imag[FSM_fft_64_stage_1_0_t1215 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1217 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010111;
    FSM_fft_64_stage_1_0_t1218 = FSM_fft_64_stage_1_0_t1217[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1219 = FSM_fft_64_stage_1_0_t1218 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1220 = FSM_fft_64_stage_1_0_t1219[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1221 = FSM_fft_64_stage_1_0_t1220[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1222 = i_data_in_imag[FSM_fft_64_stage_1_0_t1221 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1223 = FSM_fft_64_stage_1_0_t1216 + FSM_fft_64_stage_1_0_t1222;
    FSM_fft_64_stage_1_0_t1224 = FSM_fft_64_stage_1_0_t1223[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1225 = FSM_fft_64_stage_1_0_t1209;
    FSM_fft_64_stage_1_0_t1225[FSM_fft_64_stage_1_0_t1212 * 32 +: 32] = FSM_fft_64_stage_1_0_t1224;
    FSM_fft_64_stage_1_0_t1226 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000010111;
    FSM_fft_64_stage_1_0_t1227 = FSM_fft_64_stage_1_0_t1226[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1228 = FSM_fft_64_stage_1_0_t1227 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1229 = FSM_fft_64_stage_1_0_t1228[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1230 = FSM_fft_64_stage_1_0_t1229[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1231 = FSM_fft_64_stage_1_0_t1225;
    FSM_fft_64_stage_1_0_t1231[FSM_fft_64_stage_1_0_t1230 * 32 +: 32] = FSM_fft_64_stage_1_0_t1216 - FSM_fft_64_stage_1_0_t1222;
    FSM_fft_64_stage_1_0_t1232 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011000;
    FSM_fft_64_stage_1_0_t1233 = FSM_fft_64_stage_1_0_t1232[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1234 = FSM_fft_64_stage_1_0_t1233[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1235 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011000;
    FSM_fft_64_stage_1_0_t1236 = FSM_fft_64_stage_1_0_t1235[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1237 = FSM_fft_64_stage_1_0_t1236[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1238 = i_data_in_imag[FSM_fft_64_stage_1_0_t1237 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1239 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011000;
    FSM_fft_64_stage_1_0_t1240 = FSM_fft_64_stage_1_0_t1239[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1241 = FSM_fft_64_stage_1_0_t1240 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1242 = FSM_fft_64_stage_1_0_t1241[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1243 = FSM_fft_64_stage_1_0_t1242[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1244 = i_data_in_imag[FSM_fft_64_stage_1_0_t1243 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1245 = FSM_fft_64_stage_1_0_t1238 + FSM_fft_64_stage_1_0_t1244;
    FSM_fft_64_stage_1_0_t1246 = FSM_fft_64_stage_1_0_t1245[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1247 = FSM_fft_64_stage_1_0_t1231;
    FSM_fft_64_stage_1_0_t1247[FSM_fft_64_stage_1_0_t1234 * 32 +: 32] = FSM_fft_64_stage_1_0_t1246;
    FSM_fft_64_stage_1_0_t1248 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011000;
    FSM_fft_64_stage_1_0_t1249 = FSM_fft_64_stage_1_0_t1248[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1250 = FSM_fft_64_stage_1_0_t1249 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1251 = FSM_fft_64_stage_1_0_t1250[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1252 = FSM_fft_64_stage_1_0_t1251[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1253 = FSM_fft_64_stage_1_0_t1247;
    FSM_fft_64_stage_1_0_t1253[FSM_fft_64_stage_1_0_t1252 * 32 +: 32] = FSM_fft_64_stage_1_0_t1238 - FSM_fft_64_stage_1_0_t1244;
    FSM_fft_64_stage_1_0_t1254 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011001;
    FSM_fft_64_stage_1_0_t1255 = FSM_fft_64_stage_1_0_t1254[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1256 = FSM_fft_64_stage_1_0_t1255[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1257 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011001;
    FSM_fft_64_stage_1_0_t1258 = FSM_fft_64_stage_1_0_t1257[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1259 = FSM_fft_64_stage_1_0_t1258[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1260 = i_data_in_imag[FSM_fft_64_stage_1_0_t1259 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1261 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011001;
    FSM_fft_64_stage_1_0_t1262 = FSM_fft_64_stage_1_0_t1261[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1263 = FSM_fft_64_stage_1_0_t1262 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1264 = FSM_fft_64_stage_1_0_t1263[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1265 = FSM_fft_64_stage_1_0_t1264[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1266 = i_data_in_imag[FSM_fft_64_stage_1_0_t1265 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1267 = FSM_fft_64_stage_1_0_t1260 + FSM_fft_64_stage_1_0_t1266;
    FSM_fft_64_stage_1_0_t1268 = FSM_fft_64_stage_1_0_t1267[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1269 = FSM_fft_64_stage_1_0_t1253;
    FSM_fft_64_stage_1_0_t1269[FSM_fft_64_stage_1_0_t1256 * 32 +: 32] = FSM_fft_64_stage_1_0_t1268;
    FSM_fft_64_stage_1_0_t1270 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011001;
    FSM_fft_64_stage_1_0_t1271 = FSM_fft_64_stage_1_0_t1270[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1272 = FSM_fft_64_stage_1_0_t1271 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1273 = FSM_fft_64_stage_1_0_t1272[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1274 = FSM_fft_64_stage_1_0_t1273[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1275 = FSM_fft_64_stage_1_0_t1269;
    FSM_fft_64_stage_1_0_t1275[FSM_fft_64_stage_1_0_t1274 * 32 +: 32] = FSM_fft_64_stage_1_0_t1260 - FSM_fft_64_stage_1_0_t1266;
    FSM_fft_64_stage_1_0_t1276 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011010;
    FSM_fft_64_stage_1_0_t1277 = FSM_fft_64_stage_1_0_t1276[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1278 = FSM_fft_64_stage_1_0_t1277[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1279 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011010;
    FSM_fft_64_stage_1_0_t1280 = FSM_fft_64_stage_1_0_t1279[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1281 = FSM_fft_64_stage_1_0_t1280[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1282 = i_data_in_imag[FSM_fft_64_stage_1_0_t1281 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1283 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011010;
    FSM_fft_64_stage_1_0_t1284 = FSM_fft_64_stage_1_0_t1283[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1285 = FSM_fft_64_stage_1_0_t1284 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1286 = FSM_fft_64_stage_1_0_t1285[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1287 = FSM_fft_64_stage_1_0_t1286[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1288 = i_data_in_imag[FSM_fft_64_stage_1_0_t1287 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1289 = FSM_fft_64_stage_1_0_t1282 + FSM_fft_64_stage_1_0_t1288;
    FSM_fft_64_stage_1_0_t1290 = FSM_fft_64_stage_1_0_t1289[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1291 = FSM_fft_64_stage_1_0_t1275;
    FSM_fft_64_stage_1_0_t1291[FSM_fft_64_stage_1_0_t1278 * 32 +: 32] = FSM_fft_64_stage_1_0_t1290;
    FSM_fft_64_stage_1_0_t1292 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011010;
    FSM_fft_64_stage_1_0_t1293 = FSM_fft_64_stage_1_0_t1292[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1294 = FSM_fft_64_stage_1_0_t1293 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1295 = FSM_fft_64_stage_1_0_t1294[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1296 = FSM_fft_64_stage_1_0_t1295[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1297 = FSM_fft_64_stage_1_0_t1291;
    FSM_fft_64_stage_1_0_t1297[FSM_fft_64_stage_1_0_t1296 * 32 +: 32] = FSM_fft_64_stage_1_0_t1282 - FSM_fft_64_stage_1_0_t1288;
    FSM_fft_64_stage_1_0_t1298 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011011;
    FSM_fft_64_stage_1_0_t1299 = FSM_fft_64_stage_1_0_t1298[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1300 = FSM_fft_64_stage_1_0_t1299[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1301 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011011;
    FSM_fft_64_stage_1_0_t1302 = FSM_fft_64_stage_1_0_t1301[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1303 = FSM_fft_64_stage_1_0_t1302[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1304 = i_data_in_imag[FSM_fft_64_stage_1_0_t1303 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1305 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011011;
    FSM_fft_64_stage_1_0_t1306 = FSM_fft_64_stage_1_0_t1305[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1307 = FSM_fft_64_stage_1_0_t1306 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1308 = FSM_fft_64_stage_1_0_t1307[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1309 = FSM_fft_64_stage_1_0_t1308[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1310 = i_data_in_imag[FSM_fft_64_stage_1_0_t1309 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1311 = FSM_fft_64_stage_1_0_t1304 + FSM_fft_64_stage_1_0_t1310;
    FSM_fft_64_stage_1_0_t1312 = FSM_fft_64_stage_1_0_t1311[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1313 = FSM_fft_64_stage_1_0_t1297;
    FSM_fft_64_stage_1_0_t1313[FSM_fft_64_stage_1_0_t1300 * 32 +: 32] = FSM_fft_64_stage_1_0_t1312;
    FSM_fft_64_stage_1_0_t1314 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011011;
    FSM_fft_64_stage_1_0_t1315 = FSM_fft_64_stage_1_0_t1314[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1316 = FSM_fft_64_stage_1_0_t1315 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1317 = FSM_fft_64_stage_1_0_t1316[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1318 = FSM_fft_64_stage_1_0_t1317[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1319 = FSM_fft_64_stage_1_0_t1313;
    FSM_fft_64_stage_1_0_t1319[FSM_fft_64_stage_1_0_t1318 * 32 +: 32] = FSM_fft_64_stage_1_0_t1304 - FSM_fft_64_stage_1_0_t1310;
    FSM_fft_64_stage_1_0_t1320 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011100;
    FSM_fft_64_stage_1_0_t1321 = FSM_fft_64_stage_1_0_t1320[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1322 = FSM_fft_64_stage_1_0_t1321[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1323 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011100;
    FSM_fft_64_stage_1_0_t1324 = FSM_fft_64_stage_1_0_t1323[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1325 = FSM_fft_64_stage_1_0_t1324[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1326 = i_data_in_imag[FSM_fft_64_stage_1_0_t1325 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1327 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011100;
    FSM_fft_64_stage_1_0_t1328 = FSM_fft_64_stage_1_0_t1327[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1329 = FSM_fft_64_stage_1_0_t1328 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1330 = FSM_fft_64_stage_1_0_t1329[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1331 = FSM_fft_64_stage_1_0_t1330[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1332 = i_data_in_imag[FSM_fft_64_stage_1_0_t1331 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1333 = FSM_fft_64_stage_1_0_t1326 + FSM_fft_64_stage_1_0_t1332;
    FSM_fft_64_stage_1_0_t1334 = FSM_fft_64_stage_1_0_t1333[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1335 = FSM_fft_64_stage_1_0_t1319;
    FSM_fft_64_stage_1_0_t1335[FSM_fft_64_stage_1_0_t1322 * 32 +: 32] = FSM_fft_64_stage_1_0_t1334;
    FSM_fft_64_stage_1_0_t1336 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011100;
    FSM_fft_64_stage_1_0_t1337 = FSM_fft_64_stage_1_0_t1336[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1338 = FSM_fft_64_stage_1_0_t1337 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1339 = FSM_fft_64_stage_1_0_t1338[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1340 = FSM_fft_64_stage_1_0_t1339[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1341 = FSM_fft_64_stage_1_0_t1335;
    FSM_fft_64_stage_1_0_t1341[FSM_fft_64_stage_1_0_t1340 * 32 +: 32] = FSM_fft_64_stage_1_0_t1326 - FSM_fft_64_stage_1_0_t1332;
    FSM_fft_64_stage_1_0_t1342 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011101;
    FSM_fft_64_stage_1_0_t1343 = FSM_fft_64_stage_1_0_t1342[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1344 = FSM_fft_64_stage_1_0_t1343[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1345 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011101;
    FSM_fft_64_stage_1_0_t1346 = FSM_fft_64_stage_1_0_t1345[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1347 = FSM_fft_64_stage_1_0_t1346[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1348 = i_data_in_imag[FSM_fft_64_stage_1_0_t1347 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1349 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011101;
    FSM_fft_64_stage_1_0_t1350 = FSM_fft_64_stage_1_0_t1349[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1351 = FSM_fft_64_stage_1_0_t1350 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1352 = FSM_fft_64_stage_1_0_t1351[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1353 = FSM_fft_64_stage_1_0_t1352[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1354 = i_data_in_imag[FSM_fft_64_stage_1_0_t1353 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1355 = FSM_fft_64_stage_1_0_t1348 + FSM_fft_64_stage_1_0_t1354;
    FSM_fft_64_stage_1_0_t1356 = FSM_fft_64_stage_1_0_t1355[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1357 = FSM_fft_64_stage_1_0_t1341;
    FSM_fft_64_stage_1_0_t1357[FSM_fft_64_stage_1_0_t1344 * 32 +: 32] = FSM_fft_64_stage_1_0_t1356;
    FSM_fft_64_stage_1_0_t1358 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011101;
    FSM_fft_64_stage_1_0_t1359 = FSM_fft_64_stage_1_0_t1358[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1360 = FSM_fft_64_stage_1_0_t1359 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1361 = FSM_fft_64_stage_1_0_t1360[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1362 = FSM_fft_64_stage_1_0_t1361[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1363 = FSM_fft_64_stage_1_0_t1357;
    FSM_fft_64_stage_1_0_t1363[FSM_fft_64_stage_1_0_t1362 * 32 +: 32] = FSM_fft_64_stage_1_0_t1348 - FSM_fft_64_stage_1_0_t1354;
    FSM_fft_64_stage_1_0_t1364 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011110;
    FSM_fft_64_stage_1_0_t1365 = FSM_fft_64_stage_1_0_t1364[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1366 = FSM_fft_64_stage_1_0_t1365[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1367 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011110;
    FSM_fft_64_stage_1_0_t1368 = FSM_fft_64_stage_1_0_t1367[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1369 = FSM_fft_64_stage_1_0_t1368[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1370 = i_data_in_imag[FSM_fft_64_stage_1_0_t1369 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1371 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011110;
    FSM_fft_64_stage_1_0_t1372 = FSM_fft_64_stage_1_0_t1371[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1373 = FSM_fft_64_stage_1_0_t1372 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1374 = FSM_fft_64_stage_1_0_t1373[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1375 = FSM_fft_64_stage_1_0_t1374[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1376 = i_data_in_imag[FSM_fft_64_stage_1_0_t1375 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1377 = FSM_fft_64_stage_1_0_t1370 + FSM_fft_64_stage_1_0_t1376;
    FSM_fft_64_stage_1_0_t1378 = FSM_fft_64_stage_1_0_t1377[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1379 = FSM_fft_64_stage_1_0_t1363;
    FSM_fft_64_stage_1_0_t1379[FSM_fft_64_stage_1_0_t1366 * 32 +: 32] = FSM_fft_64_stage_1_0_t1378;
    FSM_fft_64_stage_1_0_t1380 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011110;
    FSM_fft_64_stage_1_0_t1381 = FSM_fft_64_stage_1_0_t1380[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1382 = FSM_fft_64_stage_1_0_t1381 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1383 = FSM_fft_64_stage_1_0_t1382[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1384 = FSM_fft_64_stage_1_0_t1383[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1385 = FSM_fft_64_stage_1_0_t1379;
    FSM_fft_64_stage_1_0_t1385[FSM_fft_64_stage_1_0_t1384 * 32 +: 32] = FSM_fft_64_stage_1_0_t1370 - FSM_fft_64_stage_1_0_t1376;
    FSM_fft_64_stage_1_0_t1386 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011111;
    FSM_fft_64_stage_1_0_t1387 = FSM_fft_64_stage_1_0_t1386[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1388 = FSM_fft_64_stage_1_0_t1387[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1389 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011111;
    FSM_fft_64_stage_1_0_t1390 = FSM_fft_64_stage_1_0_t1389[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1391 = FSM_fft_64_stage_1_0_t1390[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1392 = i_data_in_imag[FSM_fft_64_stage_1_0_t1391 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1393 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011111;
    FSM_fft_64_stage_1_0_t1394 = FSM_fft_64_stage_1_0_t1393[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1395 = FSM_fft_64_stage_1_0_t1394 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1396 = FSM_fft_64_stage_1_0_t1395[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1397 = FSM_fft_64_stage_1_0_t1396[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1398 = i_data_in_imag[FSM_fft_64_stage_1_0_t1397 * 32 +: 32];
    FSM_fft_64_stage_1_0_t1399 = FSM_fft_64_stage_1_0_t1392 + FSM_fft_64_stage_1_0_t1398;
    FSM_fft_64_stage_1_0_t1400 = FSM_fft_64_stage_1_0_t1399[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1401 = FSM_fft_64_stage_1_0_t1385;
    FSM_fft_64_stage_1_0_t1401[FSM_fft_64_stage_1_0_t1388 * 32 +: 32] = FSM_fft_64_stage_1_0_t1400;
    FSM_fft_64_stage_1_0_t1402 = 32'b00000000000000000000000000000010 * 32'b00000000000000000000000000011111;
    FSM_fft_64_stage_1_0_t1403 = FSM_fft_64_stage_1_0_t1402[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1404 = FSM_fft_64_stage_1_0_t1403 + 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_1_0_t1405 = FSM_fft_64_stage_1_0_t1404[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_1_0_t1406 = FSM_fft_64_stage_1_0_t1405[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_1_0_t1407 = FSM_fft_64_stage_1_0_t1401;
    FSM_fft_64_stage_1_0_t1407[FSM_fft_64_stage_1_0_t1406 * 32 +: 32] = FSM_fft_64_stage_1_0_t1392 - FSM_fft_64_stage_1_0_t1398;
end

assign FSM_fft_64_stage_1_0_in_ready = 1'b1;

always @(posedge clk) begin
    FSM_fft_64_stage_1_0_st_dummy_reg <= FSM_fft_64_stage_1_0_st_dummy_reg;
    if (rst) begin
        FSM_fft_64_stage_1_0_st_dummy_reg <= 32'b0;
    end
end
/* End submodules of fft_64_stage_1 */
/* End module fft_64_stage_1 */
endgenerate
endmodule
