`timescale 1ns / 1ps

module fft_64_stage_6_inner
(
    input wire clk,
    input wire rst,
    input wire [2048-1:0] i_data_in_real,
    input wire [2048-1:0] i_data_in_imag,
    input wire i_valid,
    output wire i_ready,
    output wire [2048-1:0] o_data_out_real,
    output wire [2048-1:0] o_data_out_imag,
    output wire o_valid,
    input wire o_ready
);

generate
/*
    Begin module fft_64_stage_6
*/
/*
    Wires declared by fft_64_stage_6
*/
wire FSM_fft_64_stage_6_0_in_ready;
wire FSM_fft_64_stage_6_0_out_valid;
/* End wires declared by fft_64_stage_6 */


/*
    Submodules of fft_64_stage_6
*/
reg [32-1:0] FSM_fft_64_stage_6_0_st_dummy_reg = 32'b0;

reg [32-1:0] FSM_fft_64_stage_6_0_t0;
reg [6-1:0] FSM_fft_64_stage_6_0_t1;
reg [32-1:0] FSM_fft_64_stage_6_0_t2;
reg [6-1:0] FSM_fft_64_stage_6_0_t3;
reg [32-1:0] FSM_fft_64_stage_6_0_t4;
reg [32-1:0] FSM_fft_64_stage_6_0_t5;
reg [6-1:0] FSM_fft_64_stage_6_0_t6;
reg [32-1:0] FSM_fft_64_stage_6_0_t7;
reg [33-1:0] FSM_fft_64_stage_6_0_t8;
reg [32-1:0] FSM_fft_64_stage_6_0_t9;
reg [2048-1:0] FSM_fft_64_stage_6_0_t10;
reg [32-1:0] FSM_fft_64_stage_6_0_t11;
reg [6-1:0] FSM_fft_64_stage_6_0_t12;
reg [32-1:0] FSM_fft_64_stage_6_0_t13;
reg [6-1:0] FSM_fft_64_stage_6_0_t14;
reg [32-1:0] FSM_fft_64_stage_6_0_t15;
reg [32-1:0] FSM_fft_64_stage_6_0_t16;
reg [6-1:0] FSM_fft_64_stage_6_0_t17;
reg [32-1:0] FSM_fft_64_stage_6_0_t18;
reg [2048-1:0] FSM_fft_64_stage_6_0_t19;
reg [32-1:0] FSM_fft_64_stage_6_0_t20;
reg [6-1:0] FSM_fft_64_stage_6_0_t21;
reg [32-1:0] FSM_fft_64_stage_6_0_t22;
reg [6-1:0] FSM_fft_64_stage_6_0_t23;
reg [32-1:0] FSM_fft_64_stage_6_0_t24;
reg [32-1:0] FSM_fft_64_stage_6_0_t25;
reg [6-1:0] FSM_fft_64_stage_6_0_t26;
reg [32-1:0] FSM_fft_64_stage_6_0_t27;
reg [33-1:0] FSM_fft_64_stage_6_0_t28;
reg [32-1:0] FSM_fft_64_stage_6_0_t29;
reg [2048-1:0] FSM_fft_64_stage_6_0_t30;
reg [32-1:0] FSM_fft_64_stage_6_0_t31;
reg [6-1:0] FSM_fft_64_stage_6_0_t32;
reg [32-1:0] FSM_fft_64_stage_6_0_t33;
reg [6-1:0] FSM_fft_64_stage_6_0_t34;
reg [32-1:0] FSM_fft_64_stage_6_0_t35;
reg [32-1:0] FSM_fft_64_stage_6_0_t36;
reg [6-1:0] FSM_fft_64_stage_6_0_t37;
reg [32-1:0] FSM_fft_64_stage_6_0_t38;
reg [2048-1:0] FSM_fft_64_stage_6_0_t39;
reg [32-1:0] FSM_fft_64_stage_6_0_t40;
reg [6-1:0] FSM_fft_64_stage_6_0_t41;
reg [32-1:0] FSM_fft_64_stage_6_0_t42;
reg [6-1:0] FSM_fft_64_stage_6_0_t43;
reg [32-1:0] FSM_fft_64_stage_6_0_t44;
reg [32-1:0] FSM_fft_64_stage_6_0_t45;
reg [6-1:0] FSM_fft_64_stage_6_0_t46;
reg [32-1:0] FSM_fft_64_stage_6_0_t47;
reg [33-1:0] FSM_fft_64_stage_6_0_t48;
reg [32-1:0] FSM_fft_64_stage_6_0_t49;
reg [2048-1:0] FSM_fft_64_stage_6_0_t50;
reg [32-1:0] FSM_fft_64_stage_6_0_t51;
reg [6-1:0] FSM_fft_64_stage_6_0_t52;
reg [32-1:0] FSM_fft_64_stage_6_0_t53;
reg [6-1:0] FSM_fft_64_stage_6_0_t54;
reg [32-1:0] FSM_fft_64_stage_6_0_t55;
reg [32-1:0] FSM_fft_64_stage_6_0_t56;
reg [6-1:0] FSM_fft_64_stage_6_0_t57;
reg [32-1:0] FSM_fft_64_stage_6_0_t58;
reg [2048-1:0] FSM_fft_64_stage_6_0_t59;
reg [32-1:0] FSM_fft_64_stage_6_0_t60;
reg [6-1:0] FSM_fft_64_stage_6_0_t61;
reg [32-1:0] FSM_fft_64_stage_6_0_t62;
reg [6-1:0] FSM_fft_64_stage_6_0_t63;
reg [32-1:0] FSM_fft_64_stage_6_0_t64;
reg [32-1:0] FSM_fft_64_stage_6_0_t65;
reg [6-1:0] FSM_fft_64_stage_6_0_t66;
reg [32-1:0] FSM_fft_64_stage_6_0_t67;
reg [33-1:0] FSM_fft_64_stage_6_0_t68;
reg [32-1:0] FSM_fft_64_stage_6_0_t69;
reg [2048-1:0] FSM_fft_64_stage_6_0_t70;
reg [32-1:0] FSM_fft_64_stage_6_0_t71;
reg [6-1:0] FSM_fft_64_stage_6_0_t72;
reg [32-1:0] FSM_fft_64_stage_6_0_t73;
reg [6-1:0] FSM_fft_64_stage_6_0_t74;
reg [32-1:0] FSM_fft_64_stage_6_0_t75;
reg [32-1:0] FSM_fft_64_stage_6_0_t76;
reg [6-1:0] FSM_fft_64_stage_6_0_t77;
reg [32-1:0] FSM_fft_64_stage_6_0_t78;
reg [2048-1:0] FSM_fft_64_stage_6_0_t79;
reg [32-1:0] FSM_fft_64_stage_6_0_t80;
reg [6-1:0] FSM_fft_64_stage_6_0_t81;
reg [32-1:0] FSM_fft_64_stage_6_0_t82;
reg [6-1:0] FSM_fft_64_stage_6_0_t83;
reg [32-1:0] FSM_fft_64_stage_6_0_t84;
reg [32-1:0] FSM_fft_64_stage_6_0_t85;
reg [6-1:0] FSM_fft_64_stage_6_0_t86;
reg [32-1:0] FSM_fft_64_stage_6_0_t87;
reg [33-1:0] FSM_fft_64_stage_6_0_t88;
reg [32-1:0] FSM_fft_64_stage_6_0_t89;
reg [2048-1:0] FSM_fft_64_stage_6_0_t90;
reg [32-1:0] FSM_fft_64_stage_6_0_t91;
reg [6-1:0] FSM_fft_64_stage_6_0_t92;
reg [32-1:0] FSM_fft_64_stage_6_0_t93;
reg [6-1:0] FSM_fft_64_stage_6_0_t94;
reg [32-1:0] FSM_fft_64_stage_6_0_t95;
reg [32-1:0] FSM_fft_64_stage_6_0_t96;
reg [6-1:0] FSM_fft_64_stage_6_0_t97;
reg [32-1:0] FSM_fft_64_stage_6_0_t98;
reg [2048-1:0] FSM_fft_64_stage_6_0_t99;
reg [32-1:0] FSM_fft_64_stage_6_0_t100;
reg [6-1:0] FSM_fft_64_stage_6_0_t101;
reg [32-1:0] FSM_fft_64_stage_6_0_t102;
reg [6-1:0] FSM_fft_64_stage_6_0_t103;
reg [32-1:0] FSM_fft_64_stage_6_0_t104;
reg [32-1:0] FSM_fft_64_stage_6_0_t105;
reg [6-1:0] FSM_fft_64_stage_6_0_t106;
reg [32-1:0] FSM_fft_64_stage_6_0_t107;
reg [33-1:0] FSM_fft_64_stage_6_0_t108;
reg [32-1:0] FSM_fft_64_stage_6_0_t109;
reg [2048-1:0] FSM_fft_64_stage_6_0_t110;
reg [32-1:0] FSM_fft_64_stage_6_0_t111;
reg [6-1:0] FSM_fft_64_stage_6_0_t112;
reg [32-1:0] FSM_fft_64_stage_6_0_t113;
reg [6-1:0] FSM_fft_64_stage_6_0_t114;
reg [32-1:0] FSM_fft_64_stage_6_0_t115;
reg [32-1:0] FSM_fft_64_stage_6_0_t116;
reg [6-1:0] FSM_fft_64_stage_6_0_t117;
reg [32-1:0] FSM_fft_64_stage_6_0_t118;
reg [2048-1:0] FSM_fft_64_stage_6_0_t119;
reg [32-1:0] FSM_fft_64_stage_6_0_t120;
reg [6-1:0] FSM_fft_64_stage_6_0_t121;
reg [32-1:0] FSM_fft_64_stage_6_0_t122;
reg [6-1:0] FSM_fft_64_stage_6_0_t123;
reg [32-1:0] FSM_fft_64_stage_6_0_t124;
reg [32-1:0] FSM_fft_64_stage_6_0_t125;
reg [6-1:0] FSM_fft_64_stage_6_0_t126;
reg [32-1:0] FSM_fft_64_stage_6_0_t127;
reg [33-1:0] FSM_fft_64_stage_6_0_t128;
reg [32-1:0] FSM_fft_64_stage_6_0_t129;
reg [2048-1:0] FSM_fft_64_stage_6_0_t130;
reg [32-1:0] FSM_fft_64_stage_6_0_t131;
reg [6-1:0] FSM_fft_64_stage_6_0_t132;
reg [32-1:0] FSM_fft_64_stage_6_0_t133;
reg [6-1:0] FSM_fft_64_stage_6_0_t134;
reg [32-1:0] FSM_fft_64_stage_6_0_t135;
reg [32-1:0] FSM_fft_64_stage_6_0_t136;
reg [6-1:0] FSM_fft_64_stage_6_0_t137;
reg [32-1:0] FSM_fft_64_stage_6_0_t138;
reg [2048-1:0] FSM_fft_64_stage_6_0_t139;
reg [32-1:0] FSM_fft_64_stage_6_0_t140;
reg [6-1:0] FSM_fft_64_stage_6_0_t141;
reg [32-1:0] FSM_fft_64_stage_6_0_t142;
reg [6-1:0] FSM_fft_64_stage_6_0_t143;
reg [32-1:0] FSM_fft_64_stage_6_0_t144;
reg [32-1:0] FSM_fft_64_stage_6_0_t145;
reg [6-1:0] FSM_fft_64_stage_6_0_t146;
reg [32-1:0] FSM_fft_64_stage_6_0_t147;
reg [33-1:0] FSM_fft_64_stage_6_0_t148;
reg [32-1:0] FSM_fft_64_stage_6_0_t149;
reg [2048-1:0] FSM_fft_64_stage_6_0_t150;
reg [32-1:0] FSM_fft_64_stage_6_0_t151;
reg [6-1:0] FSM_fft_64_stage_6_0_t152;
reg [32-1:0] FSM_fft_64_stage_6_0_t153;
reg [6-1:0] FSM_fft_64_stage_6_0_t154;
reg [32-1:0] FSM_fft_64_stage_6_0_t155;
reg [32-1:0] FSM_fft_64_stage_6_0_t156;
reg [6-1:0] FSM_fft_64_stage_6_0_t157;
reg [32-1:0] FSM_fft_64_stage_6_0_t158;
reg [2048-1:0] FSM_fft_64_stage_6_0_t159;
reg [32-1:0] FSM_fft_64_stage_6_0_t160;
reg [6-1:0] FSM_fft_64_stage_6_0_t161;
reg [32-1:0] FSM_fft_64_stage_6_0_t162;
reg [6-1:0] FSM_fft_64_stage_6_0_t163;
reg [32-1:0] FSM_fft_64_stage_6_0_t164;
reg [32-1:0] FSM_fft_64_stage_6_0_t165;
reg [6-1:0] FSM_fft_64_stage_6_0_t166;
reg [32-1:0] FSM_fft_64_stage_6_0_t167;
reg [33-1:0] FSM_fft_64_stage_6_0_t168;
reg [32-1:0] FSM_fft_64_stage_6_0_t169;
reg [2048-1:0] FSM_fft_64_stage_6_0_t170;
reg [32-1:0] FSM_fft_64_stage_6_0_t171;
reg [6-1:0] FSM_fft_64_stage_6_0_t172;
reg [32-1:0] FSM_fft_64_stage_6_0_t173;
reg [6-1:0] FSM_fft_64_stage_6_0_t174;
reg [32-1:0] FSM_fft_64_stage_6_0_t175;
reg [32-1:0] FSM_fft_64_stage_6_0_t176;
reg [6-1:0] FSM_fft_64_stage_6_0_t177;
reg [32-1:0] FSM_fft_64_stage_6_0_t178;
reg [2048-1:0] FSM_fft_64_stage_6_0_t179;
reg [32-1:0] FSM_fft_64_stage_6_0_t180;
reg [6-1:0] FSM_fft_64_stage_6_0_t181;
reg [32-1:0] FSM_fft_64_stage_6_0_t182;
reg [6-1:0] FSM_fft_64_stage_6_0_t183;
reg [32-1:0] FSM_fft_64_stage_6_0_t184;
reg [32-1:0] FSM_fft_64_stage_6_0_t185;
reg [6-1:0] FSM_fft_64_stage_6_0_t186;
reg [32-1:0] FSM_fft_64_stage_6_0_t187;
reg [33-1:0] FSM_fft_64_stage_6_0_t188;
reg [32-1:0] FSM_fft_64_stage_6_0_t189;
reg [2048-1:0] FSM_fft_64_stage_6_0_t190;
reg [32-1:0] FSM_fft_64_stage_6_0_t191;
reg [6-1:0] FSM_fft_64_stage_6_0_t192;
reg [32-1:0] FSM_fft_64_stage_6_0_t193;
reg [6-1:0] FSM_fft_64_stage_6_0_t194;
reg [32-1:0] FSM_fft_64_stage_6_0_t195;
reg [32-1:0] FSM_fft_64_stage_6_0_t196;
reg [6-1:0] FSM_fft_64_stage_6_0_t197;
reg [32-1:0] FSM_fft_64_stage_6_0_t198;
reg [2048-1:0] FSM_fft_64_stage_6_0_t199;
reg [32-1:0] FSM_fft_64_stage_6_0_t200;
reg [6-1:0] FSM_fft_64_stage_6_0_t201;
reg [32-1:0] FSM_fft_64_stage_6_0_t202;
reg [6-1:0] FSM_fft_64_stage_6_0_t203;
reg [32-1:0] FSM_fft_64_stage_6_0_t204;
reg [32-1:0] FSM_fft_64_stage_6_0_t205;
reg [6-1:0] FSM_fft_64_stage_6_0_t206;
reg [32-1:0] FSM_fft_64_stage_6_0_t207;
reg [33-1:0] FSM_fft_64_stage_6_0_t208;
reg [32-1:0] FSM_fft_64_stage_6_0_t209;
reg [2048-1:0] FSM_fft_64_stage_6_0_t210;
reg [32-1:0] FSM_fft_64_stage_6_0_t211;
reg [6-1:0] FSM_fft_64_stage_6_0_t212;
reg [32-1:0] FSM_fft_64_stage_6_0_t213;
reg [6-1:0] FSM_fft_64_stage_6_0_t214;
reg [32-1:0] FSM_fft_64_stage_6_0_t215;
reg [32-1:0] FSM_fft_64_stage_6_0_t216;
reg [6-1:0] FSM_fft_64_stage_6_0_t217;
reg [32-1:0] FSM_fft_64_stage_6_0_t218;
reg [2048-1:0] FSM_fft_64_stage_6_0_t219;
reg [32-1:0] FSM_fft_64_stage_6_0_t220;
reg [6-1:0] FSM_fft_64_stage_6_0_t221;
reg [32-1:0] FSM_fft_64_stage_6_0_t222;
reg [6-1:0] FSM_fft_64_stage_6_0_t223;
reg [32-1:0] FSM_fft_64_stage_6_0_t224;
reg [32-1:0] FSM_fft_64_stage_6_0_t225;
reg [6-1:0] FSM_fft_64_stage_6_0_t226;
reg [32-1:0] FSM_fft_64_stage_6_0_t227;
reg [33-1:0] FSM_fft_64_stage_6_0_t228;
reg [32-1:0] FSM_fft_64_stage_6_0_t229;
reg [2048-1:0] FSM_fft_64_stage_6_0_t230;
reg [32-1:0] FSM_fft_64_stage_6_0_t231;
reg [6-1:0] FSM_fft_64_stage_6_0_t232;
reg [32-1:0] FSM_fft_64_stage_6_0_t233;
reg [6-1:0] FSM_fft_64_stage_6_0_t234;
reg [32-1:0] FSM_fft_64_stage_6_0_t235;
reg [32-1:0] FSM_fft_64_stage_6_0_t236;
reg [6-1:0] FSM_fft_64_stage_6_0_t237;
reg [32-1:0] FSM_fft_64_stage_6_0_t238;
reg [2048-1:0] FSM_fft_64_stage_6_0_t239;
reg [32-1:0] FSM_fft_64_stage_6_0_t240;
reg [6-1:0] FSM_fft_64_stage_6_0_t241;
reg [32-1:0] FSM_fft_64_stage_6_0_t242;
reg [6-1:0] FSM_fft_64_stage_6_0_t243;
reg [32-1:0] FSM_fft_64_stage_6_0_t244;
reg [32-1:0] FSM_fft_64_stage_6_0_t245;
reg [6-1:0] FSM_fft_64_stage_6_0_t246;
reg [32-1:0] FSM_fft_64_stage_6_0_t247;
reg [33-1:0] FSM_fft_64_stage_6_0_t248;
reg [32-1:0] FSM_fft_64_stage_6_0_t249;
reg [2048-1:0] FSM_fft_64_stage_6_0_t250;
reg [32-1:0] FSM_fft_64_stage_6_0_t251;
reg [6-1:0] FSM_fft_64_stage_6_0_t252;
reg [32-1:0] FSM_fft_64_stage_6_0_t253;
reg [6-1:0] FSM_fft_64_stage_6_0_t254;
reg [32-1:0] FSM_fft_64_stage_6_0_t255;
reg [32-1:0] FSM_fft_64_stage_6_0_t256;
reg [6-1:0] FSM_fft_64_stage_6_0_t257;
reg [32-1:0] FSM_fft_64_stage_6_0_t258;
reg [2048-1:0] FSM_fft_64_stage_6_0_t259;
reg [32-1:0] FSM_fft_64_stage_6_0_t260;
reg [6-1:0] FSM_fft_64_stage_6_0_t261;
reg [32-1:0] FSM_fft_64_stage_6_0_t262;
reg [6-1:0] FSM_fft_64_stage_6_0_t263;
reg [32-1:0] FSM_fft_64_stage_6_0_t264;
reg [32-1:0] FSM_fft_64_stage_6_0_t265;
reg [6-1:0] FSM_fft_64_stage_6_0_t266;
reg [32-1:0] FSM_fft_64_stage_6_0_t267;
reg [33-1:0] FSM_fft_64_stage_6_0_t268;
reg [32-1:0] FSM_fft_64_stage_6_0_t269;
reg [2048-1:0] FSM_fft_64_stage_6_0_t270;
reg [32-1:0] FSM_fft_64_stage_6_0_t271;
reg [6-1:0] FSM_fft_64_stage_6_0_t272;
reg [32-1:0] FSM_fft_64_stage_6_0_t273;
reg [6-1:0] FSM_fft_64_stage_6_0_t274;
reg [32-1:0] FSM_fft_64_stage_6_0_t275;
reg [32-1:0] FSM_fft_64_stage_6_0_t276;
reg [6-1:0] FSM_fft_64_stage_6_0_t277;
reg [32-1:0] FSM_fft_64_stage_6_0_t278;
reg [2048-1:0] FSM_fft_64_stage_6_0_t279;
reg [32-1:0] FSM_fft_64_stage_6_0_t280;
reg [6-1:0] FSM_fft_64_stage_6_0_t281;
reg [32-1:0] FSM_fft_64_stage_6_0_t282;
reg [6-1:0] FSM_fft_64_stage_6_0_t283;
reg [32-1:0] FSM_fft_64_stage_6_0_t284;
reg [32-1:0] FSM_fft_64_stage_6_0_t285;
reg [6-1:0] FSM_fft_64_stage_6_0_t286;
reg [32-1:0] FSM_fft_64_stage_6_0_t287;
reg [33-1:0] FSM_fft_64_stage_6_0_t288;
reg [32-1:0] FSM_fft_64_stage_6_0_t289;
reg [2048-1:0] FSM_fft_64_stage_6_0_t290;
reg [32-1:0] FSM_fft_64_stage_6_0_t291;
reg [6-1:0] FSM_fft_64_stage_6_0_t292;
reg [32-1:0] FSM_fft_64_stage_6_0_t293;
reg [6-1:0] FSM_fft_64_stage_6_0_t294;
reg [32-1:0] FSM_fft_64_stage_6_0_t295;
reg [32-1:0] FSM_fft_64_stage_6_0_t296;
reg [6-1:0] FSM_fft_64_stage_6_0_t297;
reg [32-1:0] FSM_fft_64_stage_6_0_t298;
reg [2048-1:0] FSM_fft_64_stage_6_0_t299;
reg [32-1:0] FSM_fft_64_stage_6_0_t300;
reg [6-1:0] FSM_fft_64_stage_6_0_t301;
reg [32-1:0] FSM_fft_64_stage_6_0_t302;
reg [6-1:0] FSM_fft_64_stage_6_0_t303;
reg [32-1:0] FSM_fft_64_stage_6_0_t304;
reg [32-1:0] FSM_fft_64_stage_6_0_t305;
reg [6-1:0] FSM_fft_64_stage_6_0_t306;
reg [32-1:0] FSM_fft_64_stage_6_0_t307;
reg [33-1:0] FSM_fft_64_stage_6_0_t308;
reg [32-1:0] FSM_fft_64_stage_6_0_t309;
reg [2048-1:0] FSM_fft_64_stage_6_0_t310;
reg [32-1:0] FSM_fft_64_stage_6_0_t311;
reg [6-1:0] FSM_fft_64_stage_6_0_t312;
reg [32-1:0] FSM_fft_64_stage_6_0_t313;
reg [6-1:0] FSM_fft_64_stage_6_0_t314;
reg [32-1:0] FSM_fft_64_stage_6_0_t315;
reg [32-1:0] FSM_fft_64_stage_6_0_t316;
reg [6-1:0] FSM_fft_64_stage_6_0_t317;
reg [32-1:0] FSM_fft_64_stage_6_0_t318;
reg [2048-1:0] FSM_fft_64_stage_6_0_t319;
reg [32-1:0] FSM_fft_64_stage_6_0_t320;
reg [6-1:0] FSM_fft_64_stage_6_0_t321;
reg [32-1:0] FSM_fft_64_stage_6_0_t322;
reg [6-1:0] FSM_fft_64_stage_6_0_t323;
reg [32-1:0] FSM_fft_64_stage_6_0_t324;
reg [32-1:0] FSM_fft_64_stage_6_0_t325;
reg [6-1:0] FSM_fft_64_stage_6_0_t326;
reg [32-1:0] FSM_fft_64_stage_6_0_t327;
reg [33-1:0] FSM_fft_64_stage_6_0_t328;
reg [32-1:0] FSM_fft_64_stage_6_0_t329;
reg [2048-1:0] FSM_fft_64_stage_6_0_t330;
reg [32-1:0] FSM_fft_64_stage_6_0_t331;
reg [6-1:0] FSM_fft_64_stage_6_0_t332;
reg [32-1:0] FSM_fft_64_stage_6_0_t333;
reg [6-1:0] FSM_fft_64_stage_6_0_t334;
reg [32-1:0] FSM_fft_64_stage_6_0_t335;
reg [32-1:0] FSM_fft_64_stage_6_0_t336;
reg [6-1:0] FSM_fft_64_stage_6_0_t337;
reg [32-1:0] FSM_fft_64_stage_6_0_t338;
reg [2048-1:0] FSM_fft_64_stage_6_0_t339;
reg [32-1:0] FSM_fft_64_stage_6_0_t340;
reg [6-1:0] FSM_fft_64_stage_6_0_t341;
reg [32-1:0] FSM_fft_64_stage_6_0_t342;
reg [6-1:0] FSM_fft_64_stage_6_0_t343;
reg [32-1:0] FSM_fft_64_stage_6_0_t344;
reg [32-1:0] FSM_fft_64_stage_6_0_t345;
reg [6-1:0] FSM_fft_64_stage_6_0_t346;
reg [32-1:0] FSM_fft_64_stage_6_0_t347;
reg [33-1:0] FSM_fft_64_stage_6_0_t348;
reg [32-1:0] FSM_fft_64_stage_6_0_t349;
reg [2048-1:0] FSM_fft_64_stage_6_0_t350;
reg [32-1:0] FSM_fft_64_stage_6_0_t351;
reg [6-1:0] FSM_fft_64_stage_6_0_t352;
reg [32-1:0] FSM_fft_64_stage_6_0_t353;
reg [6-1:0] FSM_fft_64_stage_6_0_t354;
reg [32-1:0] FSM_fft_64_stage_6_0_t355;
reg [32-1:0] FSM_fft_64_stage_6_0_t356;
reg [6-1:0] FSM_fft_64_stage_6_0_t357;
reg [32-1:0] FSM_fft_64_stage_6_0_t358;
reg [2048-1:0] FSM_fft_64_stage_6_0_t359;
reg [32-1:0] FSM_fft_64_stage_6_0_t360;
reg [6-1:0] FSM_fft_64_stage_6_0_t361;
reg [32-1:0] FSM_fft_64_stage_6_0_t362;
reg [6-1:0] FSM_fft_64_stage_6_0_t363;
reg [32-1:0] FSM_fft_64_stage_6_0_t364;
reg [32-1:0] FSM_fft_64_stage_6_0_t365;
reg [6-1:0] FSM_fft_64_stage_6_0_t366;
reg [32-1:0] FSM_fft_64_stage_6_0_t367;
reg [33-1:0] FSM_fft_64_stage_6_0_t368;
reg [32-1:0] FSM_fft_64_stage_6_0_t369;
reg [2048-1:0] FSM_fft_64_stage_6_0_t370;
reg [32-1:0] FSM_fft_64_stage_6_0_t371;
reg [6-1:0] FSM_fft_64_stage_6_0_t372;
reg [32-1:0] FSM_fft_64_stage_6_0_t373;
reg [6-1:0] FSM_fft_64_stage_6_0_t374;
reg [32-1:0] FSM_fft_64_stage_6_0_t375;
reg [32-1:0] FSM_fft_64_stage_6_0_t376;
reg [6-1:0] FSM_fft_64_stage_6_0_t377;
reg [32-1:0] FSM_fft_64_stage_6_0_t378;
reg [2048-1:0] FSM_fft_64_stage_6_0_t379;
reg [32-1:0] FSM_fft_64_stage_6_0_t380;
reg [6-1:0] FSM_fft_64_stage_6_0_t381;
reg [32-1:0] FSM_fft_64_stage_6_0_t382;
reg [6-1:0] FSM_fft_64_stage_6_0_t383;
reg [32-1:0] FSM_fft_64_stage_6_0_t384;
reg [32-1:0] FSM_fft_64_stage_6_0_t385;
reg [6-1:0] FSM_fft_64_stage_6_0_t386;
reg [32-1:0] FSM_fft_64_stage_6_0_t387;
reg [33-1:0] FSM_fft_64_stage_6_0_t388;
reg [32-1:0] FSM_fft_64_stage_6_0_t389;
reg [2048-1:0] FSM_fft_64_stage_6_0_t390;
reg [32-1:0] FSM_fft_64_stage_6_0_t391;
reg [6-1:0] FSM_fft_64_stage_6_0_t392;
reg [32-1:0] FSM_fft_64_stage_6_0_t393;
reg [6-1:0] FSM_fft_64_stage_6_0_t394;
reg [32-1:0] FSM_fft_64_stage_6_0_t395;
reg [32-1:0] FSM_fft_64_stage_6_0_t396;
reg [6-1:0] FSM_fft_64_stage_6_0_t397;
reg [32-1:0] FSM_fft_64_stage_6_0_t398;
reg [2048-1:0] FSM_fft_64_stage_6_0_t399;
reg [32-1:0] FSM_fft_64_stage_6_0_t400;
reg [6-1:0] FSM_fft_64_stage_6_0_t401;
reg [32-1:0] FSM_fft_64_stage_6_0_t402;
reg [6-1:0] FSM_fft_64_stage_6_0_t403;
reg [32-1:0] FSM_fft_64_stage_6_0_t404;
reg [32-1:0] FSM_fft_64_stage_6_0_t405;
reg [6-1:0] FSM_fft_64_stage_6_0_t406;
reg [32-1:0] FSM_fft_64_stage_6_0_t407;
reg [33-1:0] FSM_fft_64_stage_6_0_t408;
reg [32-1:0] FSM_fft_64_stage_6_0_t409;
reg [2048-1:0] FSM_fft_64_stage_6_0_t410;
reg [32-1:0] FSM_fft_64_stage_6_0_t411;
reg [6-1:0] FSM_fft_64_stage_6_0_t412;
reg [32-1:0] FSM_fft_64_stage_6_0_t413;
reg [6-1:0] FSM_fft_64_stage_6_0_t414;
reg [32-1:0] FSM_fft_64_stage_6_0_t415;
reg [32-1:0] FSM_fft_64_stage_6_0_t416;
reg [6-1:0] FSM_fft_64_stage_6_0_t417;
reg [32-1:0] FSM_fft_64_stage_6_0_t418;
reg [2048-1:0] FSM_fft_64_stage_6_0_t419;
reg [32-1:0] FSM_fft_64_stage_6_0_t420;
reg [6-1:0] FSM_fft_64_stage_6_0_t421;
reg [32-1:0] FSM_fft_64_stage_6_0_t422;
reg [6-1:0] FSM_fft_64_stage_6_0_t423;
reg [32-1:0] FSM_fft_64_stage_6_0_t424;
reg [32-1:0] FSM_fft_64_stage_6_0_t425;
reg [6-1:0] FSM_fft_64_stage_6_0_t426;
reg [32-1:0] FSM_fft_64_stage_6_0_t427;
reg [33-1:0] FSM_fft_64_stage_6_0_t428;
reg [32-1:0] FSM_fft_64_stage_6_0_t429;
reg [2048-1:0] FSM_fft_64_stage_6_0_t430;
reg [32-1:0] FSM_fft_64_stage_6_0_t431;
reg [6-1:0] FSM_fft_64_stage_6_0_t432;
reg [32-1:0] FSM_fft_64_stage_6_0_t433;
reg [6-1:0] FSM_fft_64_stage_6_0_t434;
reg [32-1:0] FSM_fft_64_stage_6_0_t435;
reg [32-1:0] FSM_fft_64_stage_6_0_t436;
reg [6-1:0] FSM_fft_64_stage_6_0_t437;
reg [32-1:0] FSM_fft_64_stage_6_0_t438;
reg [2048-1:0] FSM_fft_64_stage_6_0_t439;
reg [32-1:0] FSM_fft_64_stage_6_0_t440;
reg [6-1:0] FSM_fft_64_stage_6_0_t441;
reg [32-1:0] FSM_fft_64_stage_6_0_t442;
reg [6-1:0] FSM_fft_64_stage_6_0_t443;
reg [32-1:0] FSM_fft_64_stage_6_0_t444;
reg [32-1:0] FSM_fft_64_stage_6_0_t445;
reg [6-1:0] FSM_fft_64_stage_6_0_t446;
reg [32-1:0] FSM_fft_64_stage_6_0_t447;
reg [33-1:0] FSM_fft_64_stage_6_0_t448;
reg [32-1:0] FSM_fft_64_stage_6_0_t449;
reg [2048-1:0] FSM_fft_64_stage_6_0_t450;
reg [32-1:0] FSM_fft_64_stage_6_0_t451;
reg [6-1:0] FSM_fft_64_stage_6_0_t452;
reg [32-1:0] FSM_fft_64_stage_6_0_t453;
reg [6-1:0] FSM_fft_64_stage_6_0_t454;
reg [32-1:0] FSM_fft_64_stage_6_0_t455;
reg [32-1:0] FSM_fft_64_stage_6_0_t456;
reg [6-1:0] FSM_fft_64_stage_6_0_t457;
reg [32-1:0] FSM_fft_64_stage_6_0_t458;
reg [2048-1:0] FSM_fft_64_stage_6_0_t459;
reg [32-1:0] FSM_fft_64_stage_6_0_t460;
reg [6-1:0] FSM_fft_64_stage_6_0_t461;
reg [32-1:0] FSM_fft_64_stage_6_0_t462;
reg [6-1:0] FSM_fft_64_stage_6_0_t463;
reg [32-1:0] FSM_fft_64_stage_6_0_t464;
reg [32-1:0] FSM_fft_64_stage_6_0_t465;
reg [6-1:0] FSM_fft_64_stage_6_0_t466;
reg [32-1:0] FSM_fft_64_stage_6_0_t467;
reg [33-1:0] FSM_fft_64_stage_6_0_t468;
reg [32-1:0] FSM_fft_64_stage_6_0_t469;
reg [2048-1:0] FSM_fft_64_stage_6_0_t470;
reg [32-1:0] FSM_fft_64_stage_6_0_t471;
reg [6-1:0] FSM_fft_64_stage_6_0_t472;
reg [32-1:0] FSM_fft_64_stage_6_0_t473;
reg [6-1:0] FSM_fft_64_stage_6_0_t474;
reg [32-1:0] FSM_fft_64_stage_6_0_t475;
reg [32-1:0] FSM_fft_64_stage_6_0_t476;
reg [6-1:0] FSM_fft_64_stage_6_0_t477;
reg [32-1:0] FSM_fft_64_stage_6_0_t478;
reg [2048-1:0] FSM_fft_64_stage_6_0_t479;
reg [32-1:0] FSM_fft_64_stage_6_0_t480;
reg [6-1:0] FSM_fft_64_stage_6_0_t481;
reg [32-1:0] FSM_fft_64_stage_6_0_t482;
reg [6-1:0] FSM_fft_64_stage_6_0_t483;
reg [32-1:0] FSM_fft_64_stage_6_0_t484;
reg [32-1:0] FSM_fft_64_stage_6_0_t485;
reg [6-1:0] FSM_fft_64_stage_6_0_t486;
reg [32-1:0] FSM_fft_64_stage_6_0_t487;
reg [33-1:0] FSM_fft_64_stage_6_0_t488;
reg [32-1:0] FSM_fft_64_stage_6_0_t489;
reg [2048-1:0] FSM_fft_64_stage_6_0_t490;
reg [32-1:0] FSM_fft_64_stage_6_0_t491;
reg [6-1:0] FSM_fft_64_stage_6_0_t492;
reg [32-1:0] FSM_fft_64_stage_6_0_t493;
reg [6-1:0] FSM_fft_64_stage_6_0_t494;
reg [32-1:0] FSM_fft_64_stage_6_0_t495;
reg [32-1:0] FSM_fft_64_stage_6_0_t496;
reg [6-1:0] FSM_fft_64_stage_6_0_t497;
reg [32-1:0] FSM_fft_64_stage_6_0_t498;
reg [2048-1:0] FSM_fft_64_stage_6_0_t499;
reg [32-1:0] FSM_fft_64_stage_6_0_t500;
reg [6-1:0] FSM_fft_64_stage_6_0_t501;
reg [32-1:0] FSM_fft_64_stage_6_0_t502;
reg [6-1:0] FSM_fft_64_stage_6_0_t503;
reg [32-1:0] FSM_fft_64_stage_6_0_t504;
reg [32-1:0] FSM_fft_64_stage_6_0_t505;
reg [6-1:0] FSM_fft_64_stage_6_0_t506;
reg [32-1:0] FSM_fft_64_stage_6_0_t507;
reg [33-1:0] FSM_fft_64_stage_6_0_t508;
reg [32-1:0] FSM_fft_64_stage_6_0_t509;
reg [2048-1:0] FSM_fft_64_stage_6_0_t510;
reg [32-1:0] FSM_fft_64_stage_6_0_t511;
reg [6-1:0] FSM_fft_64_stage_6_0_t512;
reg [32-1:0] FSM_fft_64_stage_6_0_t513;
reg [6-1:0] FSM_fft_64_stage_6_0_t514;
reg [32-1:0] FSM_fft_64_stage_6_0_t515;
reg [32-1:0] FSM_fft_64_stage_6_0_t516;
reg [6-1:0] FSM_fft_64_stage_6_0_t517;
reg [32-1:0] FSM_fft_64_stage_6_0_t518;
reg [2048-1:0] FSM_fft_64_stage_6_0_t519;
reg [32-1:0] FSM_fft_64_stage_6_0_t520;
reg [6-1:0] FSM_fft_64_stage_6_0_t521;
reg [32-1:0] FSM_fft_64_stage_6_0_t522;
reg [6-1:0] FSM_fft_64_stage_6_0_t523;
reg [32-1:0] FSM_fft_64_stage_6_0_t524;
reg [32-1:0] FSM_fft_64_stage_6_0_t525;
reg [6-1:0] FSM_fft_64_stage_6_0_t526;
reg [32-1:0] FSM_fft_64_stage_6_0_t527;
reg [33-1:0] FSM_fft_64_stage_6_0_t528;
reg [32-1:0] FSM_fft_64_stage_6_0_t529;
reg [2048-1:0] FSM_fft_64_stage_6_0_t530;
reg [32-1:0] FSM_fft_64_stage_6_0_t531;
reg [6-1:0] FSM_fft_64_stage_6_0_t532;
reg [32-1:0] FSM_fft_64_stage_6_0_t533;
reg [6-1:0] FSM_fft_64_stage_6_0_t534;
reg [32-1:0] FSM_fft_64_stage_6_0_t535;
reg [32-1:0] FSM_fft_64_stage_6_0_t536;
reg [6-1:0] FSM_fft_64_stage_6_0_t537;
reg [32-1:0] FSM_fft_64_stage_6_0_t538;
reg [2048-1:0] FSM_fft_64_stage_6_0_t539;
reg [32-1:0] FSM_fft_64_stage_6_0_t540;
reg [6-1:0] FSM_fft_64_stage_6_0_t541;
reg [32-1:0] FSM_fft_64_stage_6_0_t542;
reg [6-1:0] FSM_fft_64_stage_6_0_t543;
reg [32-1:0] FSM_fft_64_stage_6_0_t544;
reg [32-1:0] FSM_fft_64_stage_6_0_t545;
reg [6-1:0] FSM_fft_64_stage_6_0_t546;
reg [32-1:0] FSM_fft_64_stage_6_0_t547;
reg [33-1:0] FSM_fft_64_stage_6_0_t548;
reg [32-1:0] FSM_fft_64_stage_6_0_t549;
reg [2048-1:0] FSM_fft_64_stage_6_0_t550;
reg [32-1:0] FSM_fft_64_stage_6_0_t551;
reg [6-1:0] FSM_fft_64_stage_6_0_t552;
reg [32-1:0] FSM_fft_64_stage_6_0_t553;
reg [6-1:0] FSM_fft_64_stage_6_0_t554;
reg [32-1:0] FSM_fft_64_stage_6_0_t555;
reg [32-1:0] FSM_fft_64_stage_6_0_t556;
reg [6-1:0] FSM_fft_64_stage_6_0_t557;
reg [32-1:0] FSM_fft_64_stage_6_0_t558;
reg [2048-1:0] FSM_fft_64_stage_6_0_t559;
reg [32-1:0] FSM_fft_64_stage_6_0_t560;
reg [6-1:0] FSM_fft_64_stage_6_0_t561;
reg [32-1:0] FSM_fft_64_stage_6_0_t562;
reg [6-1:0] FSM_fft_64_stage_6_0_t563;
reg [32-1:0] FSM_fft_64_stage_6_0_t564;
reg [32-1:0] FSM_fft_64_stage_6_0_t565;
reg [6-1:0] FSM_fft_64_stage_6_0_t566;
reg [32-1:0] FSM_fft_64_stage_6_0_t567;
reg [33-1:0] FSM_fft_64_stage_6_0_t568;
reg [32-1:0] FSM_fft_64_stage_6_0_t569;
reg [2048-1:0] FSM_fft_64_stage_6_0_t570;
reg [32-1:0] FSM_fft_64_stage_6_0_t571;
reg [6-1:0] FSM_fft_64_stage_6_0_t572;
reg [32-1:0] FSM_fft_64_stage_6_0_t573;
reg [6-1:0] FSM_fft_64_stage_6_0_t574;
reg [32-1:0] FSM_fft_64_stage_6_0_t575;
reg [32-1:0] FSM_fft_64_stage_6_0_t576;
reg [6-1:0] FSM_fft_64_stage_6_0_t577;
reg [32-1:0] FSM_fft_64_stage_6_0_t578;
reg [2048-1:0] FSM_fft_64_stage_6_0_t579;
reg [32-1:0] FSM_fft_64_stage_6_0_t580;
reg [6-1:0] FSM_fft_64_stage_6_0_t581;
reg [32-1:0] FSM_fft_64_stage_6_0_t582;
reg [6-1:0] FSM_fft_64_stage_6_0_t583;
reg [32-1:0] FSM_fft_64_stage_6_0_t584;
reg [32-1:0] FSM_fft_64_stage_6_0_t585;
reg [6-1:0] FSM_fft_64_stage_6_0_t586;
reg [32-1:0] FSM_fft_64_stage_6_0_t587;
reg [33-1:0] FSM_fft_64_stage_6_0_t588;
reg [32-1:0] FSM_fft_64_stage_6_0_t589;
reg [2048-1:0] FSM_fft_64_stage_6_0_t590;
reg [32-1:0] FSM_fft_64_stage_6_0_t591;
reg [6-1:0] FSM_fft_64_stage_6_0_t592;
reg [32-1:0] FSM_fft_64_stage_6_0_t593;
reg [6-1:0] FSM_fft_64_stage_6_0_t594;
reg [32-1:0] FSM_fft_64_stage_6_0_t595;
reg [32-1:0] FSM_fft_64_stage_6_0_t596;
reg [6-1:0] FSM_fft_64_stage_6_0_t597;
reg [32-1:0] FSM_fft_64_stage_6_0_t598;
reg [2048-1:0] FSM_fft_64_stage_6_0_t599;
reg [32-1:0] FSM_fft_64_stage_6_0_t600;
reg [6-1:0] FSM_fft_64_stage_6_0_t601;
reg [32-1:0] FSM_fft_64_stage_6_0_t602;
reg [6-1:0] FSM_fft_64_stage_6_0_t603;
reg [32-1:0] FSM_fft_64_stage_6_0_t604;
reg [32-1:0] FSM_fft_64_stage_6_0_t605;
reg [6-1:0] FSM_fft_64_stage_6_0_t606;
reg [32-1:0] FSM_fft_64_stage_6_0_t607;
reg [33-1:0] FSM_fft_64_stage_6_0_t608;
reg [32-1:0] FSM_fft_64_stage_6_0_t609;
reg [2048-1:0] FSM_fft_64_stage_6_0_t610;
reg [32-1:0] FSM_fft_64_stage_6_0_t611;
reg [6-1:0] FSM_fft_64_stage_6_0_t612;
reg [32-1:0] FSM_fft_64_stage_6_0_t613;
reg [6-1:0] FSM_fft_64_stage_6_0_t614;
reg [32-1:0] FSM_fft_64_stage_6_0_t615;
reg [32-1:0] FSM_fft_64_stage_6_0_t616;
reg [6-1:0] FSM_fft_64_stage_6_0_t617;
reg [32-1:0] FSM_fft_64_stage_6_0_t618;
reg [2048-1:0] FSM_fft_64_stage_6_0_t619;
reg [32-1:0] FSM_fft_64_stage_6_0_t620;
reg [6-1:0] FSM_fft_64_stage_6_0_t621;
reg [32-1:0] FSM_fft_64_stage_6_0_t622;
reg [6-1:0] FSM_fft_64_stage_6_0_t623;
reg [32-1:0] FSM_fft_64_stage_6_0_t624;
reg [32-1:0] FSM_fft_64_stage_6_0_t625;
reg [6-1:0] FSM_fft_64_stage_6_0_t626;
reg [32-1:0] FSM_fft_64_stage_6_0_t627;
reg [33-1:0] FSM_fft_64_stage_6_0_t628;
reg [32-1:0] FSM_fft_64_stage_6_0_t629;
reg [2048-1:0] FSM_fft_64_stage_6_0_t630;
reg [32-1:0] FSM_fft_64_stage_6_0_t631;
reg [6-1:0] FSM_fft_64_stage_6_0_t632;
reg [32-1:0] FSM_fft_64_stage_6_0_t633;
reg [6-1:0] FSM_fft_64_stage_6_0_t634;
reg [32-1:0] FSM_fft_64_stage_6_0_t635;
reg [32-1:0] FSM_fft_64_stage_6_0_t636;
reg [6-1:0] FSM_fft_64_stage_6_0_t637;
reg [32-1:0] FSM_fft_64_stage_6_0_t638;
reg [2048-1:0] FSM_fft_64_stage_6_0_t639;
reg [32-1:0] FSM_fft_64_stage_6_0_t640;
reg [6-1:0] FSM_fft_64_stage_6_0_t641;
reg [32-1:0] FSM_fft_64_stage_6_0_t642;
reg [6-1:0] FSM_fft_64_stage_6_0_t643;
reg [32-1:0] FSM_fft_64_stage_6_0_t644;
reg [32-1:0] FSM_fft_64_stage_6_0_t645;
reg [6-1:0] FSM_fft_64_stage_6_0_t646;
reg [32-1:0] FSM_fft_64_stage_6_0_t647;
reg [33-1:0] FSM_fft_64_stage_6_0_t648;
reg [32-1:0] FSM_fft_64_stage_6_0_t649;
reg [2048-1:0] FSM_fft_64_stage_6_0_t650;
reg [32-1:0] FSM_fft_64_stage_6_0_t651;
reg [6-1:0] FSM_fft_64_stage_6_0_t652;
reg [32-1:0] FSM_fft_64_stage_6_0_t653;
reg [6-1:0] FSM_fft_64_stage_6_0_t654;
reg [32-1:0] FSM_fft_64_stage_6_0_t655;
reg [32-1:0] FSM_fft_64_stage_6_0_t656;
reg [6-1:0] FSM_fft_64_stage_6_0_t657;
reg [32-1:0] FSM_fft_64_stage_6_0_t658;
reg [2048-1:0] FSM_fft_64_stage_6_0_t659;
reg [32-1:0] FSM_fft_64_stage_6_0_t660;
reg [6-1:0] FSM_fft_64_stage_6_0_t661;
reg [32-1:0] FSM_fft_64_stage_6_0_t662;
reg [6-1:0] FSM_fft_64_stage_6_0_t663;
reg [32-1:0] FSM_fft_64_stage_6_0_t664;
reg [32-1:0] FSM_fft_64_stage_6_0_t665;
reg [6-1:0] FSM_fft_64_stage_6_0_t666;
reg [32-1:0] FSM_fft_64_stage_6_0_t667;
reg [33-1:0] FSM_fft_64_stage_6_0_t668;
reg [32-1:0] FSM_fft_64_stage_6_0_t669;
reg [2048-1:0] FSM_fft_64_stage_6_0_t670;
reg [32-1:0] FSM_fft_64_stage_6_0_t671;
reg [6-1:0] FSM_fft_64_stage_6_0_t672;
reg [32-1:0] FSM_fft_64_stage_6_0_t673;
reg [6-1:0] FSM_fft_64_stage_6_0_t674;
reg [32-1:0] FSM_fft_64_stage_6_0_t675;
reg [32-1:0] FSM_fft_64_stage_6_0_t676;
reg [6-1:0] FSM_fft_64_stage_6_0_t677;
reg [32-1:0] FSM_fft_64_stage_6_0_t678;
reg [2048-1:0] FSM_fft_64_stage_6_0_t679;
reg [32-1:0] FSM_fft_64_stage_6_0_t680;
reg [6-1:0] FSM_fft_64_stage_6_0_t681;
reg [32-1:0] FSM_fft_64_stage_6_0_t682;
reg [6-1:0] FSM_fft_64_stage_6_0_t683;
reg [32-1:0] FSM_fft_64_stage_6_0_t684;
reg [32-1:0] FSM_fft_64_stage_6_0_t685;
reg [6-1:0] FSM_fft_64_stage_6_0_t686;
reg [32-1:0] FSM_fft_64_stage_6_0_t687;
reg [33-1:0] FSM_fft_64_stage_6_0_t688;
reg [32-1:0] FSM_fft_64_stage_6_0_t689;
reg [2048-1:0] FSM_fft_64_stage_6_0_t690;
reg [32-1:0] FSM_fft_64_stage_6_0_t691;
reg [6-1:0] FSM_fft_64_stage_6_0_t692;
reg [32-1:0] FSM_fft_64_stage_6_0_t693;
reg [6-1:0] FSM_fft_64_stage_6_0_t694;
reg [32-1:0] FSM_fft_64_stage_6_0_t695;
reg [32-1:0] FSM_fft_64_stage_6_0_t696;
reg [6-1:0] FSM_fft_64_stage_6_0_t697;
reg [32-1:0] FSM_fft_64_stage_6_0_t698;
reg [2048-1:0] FSM_fft_64_stage_6_0_t699;
reg [32-1:0] FSM_fft_64_stage_6_0_t700;
reg [6-1:0] FSM_fft_64_stage_6_0_t701;
reg [32-1:0] FSM_fft_64_stage_6_0_t702;
reg [6-1:0] FSM_fft_64_stage_6_0_t703;
reg [32-1:0] FSM_fft_64_stage_6_0_t704;
reg [32-1:0] FSM_fft_64_stage_6_0_t705;
reg [6-1:0] FSM_fft_64_stage_6_0_t706;
reg [32-1:0] FSM_fft_64_stage_6_0_t707;
reg [33-1:0] FSM_fft_64_stage_6_0_t708;
reg [32-1:0] FSM_fft_64_stage_6_0_t709;
reg [2048-1:0] FSM_fft_64_stage_6_0_t710;
reg [32-1:0] FSM_fft_64_stage_6_0_t711;
reg [6-1:0] FSM_fft_64_stage_6_0_t712;
reg [32-1:0] FSM_fft_64_stage_6_0_t713;
reg [6-1:0] FSM_fft_64_stage_6_0_t714;
reg [32-1:0] FSM_fft_64_stage_6_0_t715;
reg [32-1:0] FSM_fft_64_stage_6_0_t716;
reg [6-1:0] FSM_fft_64_stage_6_0_t717;
reg [32-1:0] FSM_fft_64_stage_6_0_t718;
reg [2048-1:0] FSM_fft_64_stage_6_0_t719;
reg [32-1:0] FSM_fft_64_stage_6_0_t720;
reg [6-1:0] FSM_fft_64_stage_6_0_t721;
reg [32-1:0] FSM_fft_64_stage_6_0_t722;
reg [6-1:0] FSM_fft_64_stage_6_0_t723;
reg [32-1:0] FSM_fft_64_stage_6_0_t724;
reg [32-1:0] FSM_fft_64_stage_6_0_t725;
reg [6-1:0] FSM_fft_64_stage_6_0_t726;
reg [32-1:0] FSM_fft_64_stage_6_0_t727;
reg [33-1:0] FSM_fft_64_stage_6_0_t728;
reg [32-1:0] FSM_fft_64_stage_6_0_t729;
reg [2048-1:0] FSM_fft_64_stage_6_0_t730;
reg [32-1:0] FSM_fft_64_stage_6_0_t731;
reg [6-1:0] FSM_fft_64_stage_6_0_t732;
reg [32-1:0] FSM_fft_64_stage_6_0_t733;
reg [6-1:0] FSM_fft_64_stage_6_0_t734;
reg [32-1:0] FSM_fft_64_stage_6_0_t735;
reg [32-1:0] FSM_fft_64_stage_6_0_t736;
reg [6-1:0] FSM_fft_64_stage_6_0_t737;
reg [32-1:0] FSM_fft_64_stage_6_0_t738;
reg [2048-1:0] FSM_fft_64_stage_6_0_t739;
reg [32-1:0] FSM_fft_64_stage_6_0_t740;
reg [6-1:0] FSM_fft_64_stage_6_0_t741;
reg [32-1:0] FSM_fft_64_stage_6_0_t742;
reg [6-1:0] FSM_fft_64_stage_6_0_t743;
reg [32-1:0] FSM_fft_64_stage_6_0_t744;
reg [32-1:0] FSM_fft_64_stage_6_0_t745;
reg [6-1:0] FSM_fft_64_stage_6_0_t746;
reg [32-1:0] FSM_fft_64_stage_6_0_t747;
reg [33-1:0] FSM_fft_64_stage_6_0_t748;
reg [32-1:0] FSM_fft_64_stage_6_0_t749;
reg [2048-1:0] FSM_fft_64_stage_6_0_t750;
reg [32-1:0] FSM_fft_64_stage_6_0_t751;
reg [6-1:0] FSM_fft_64_stage_6_0_t752;
reg [32-1:0] FSM_fft_64_stage_6_0_t753;
reg [6-1:0] FSM_fft_64_stage_6_0_t754;
reg [32-1:0] FSM_fft_64_stage_6_0_t755;
reg [32-1:0] FSM_fft_64_stage_6_0_t756;
reg [6-1:0] FSM_fft_64_stage_6_0_t757;
reg [32-1:0] FSM_fft_64_stage_6_0_t758;
reg [2048-1:0] FSM_fft_64_stage_6_0_t759;
reg [32-1:0] FSM_fft_64_stage_6_0_t760;
reg [6-1:0] FSM_fft_64_stage_6_0_t761;
reg [32-1:0] FSM_fft_64_stage_6_0_t762;
reg [6-1:0] FSM_fft_64_stage_6_0_t763;
reg [32-1:0] FSM_fft_64_stage_6_0_t764;
reg [32-1:0] FSM_fft_64_stage_6_0_t765;
reg [6-1:0] FSM_fft_64_stage_6_0_t766;
reg [32-1:0] FSM_fft_64_stage_6_0_t767;
reg [33-1:0] FSM_fft_64_stage_6_0_t768;
reg [32-1:0] FSM_fft_64_stage_6_0_t769;
reg [2048-1:0] FSM_fft_64_stage_6_0_t770;
reg [32-1:0] FSM_fft_64_stage_6_0_t771;
reg [6-1:0] FSM_fft_64_stage_6_0_t772;
reg [32-1:0] FSM_fft_64_stage_6_0_t773;
reg [6-1:0] FSM_fft_64_stage_6_0_t774;
reg [32-1:0] FSM_fft_64_stage_6_0_t775;
reg [32-1:0] FSM_fft_64_stage_6_0_t776;
reg [6-1:0] FSM_fft_64_stage_6_0_t777;
reg [32-1:0] FSM_fft_64_stage_6_0_t778;
reg [2048-1:0] FSM_fft_64_stage_6_0_t779;
reg [32-1:0] FSM_fft_64_stage_6_0_t780;
reg [6-1:0] FSM_fft_64_stage_6_0_t781;
reg [32-1:0] FSM_fft_64_stage_6_0_t782;
reg [6-1:0] FSM_fft_64_stage_6_0_t783;
reg [32-1:0] FSM_fft_64_stage_6_0_t784;
reg [32-1:0] FSM_fft_64_stage_6_0_t785;
reg [6-1:0] FSM_fft_64_stage_6_0_t786;
reg [32-1:0] FSM_fft_64_stage_6_0_t787;
reg [33-1:0] FSM_fft_64_stage_6_0_t788;
reg [32-1:0] FSM_fft_64_stage_6_0_t789;
reg [2048-1:0] FSM_fft_64_stage_6_0_t790;
reg [32-1:0] FSM_fft_64_stage_6_0_t791;
reg [6-1:0] FSM_fft_64_stage_6_0_t792;
reg [32-1:0] FSM_fft_64_stage_6_0_t793;
reg [6-1:0] FSM_fft_64_stage_6_0_t794;
reg [32-1:0] FSM_fft_64_stage_6_0_t795;
reg [32-1:0] FSM_fft_64_stage_6_0_t796;
reg [6-1:0] FSM_fft_64_stage_6_0_t797;
reg [32-1:0] FSM_fft_64_stage_6_0_t798;
reg [2048-1:0] FSM_fft_64_stage_6_0_t799;
reg [32-1:0] FSM_fft_64_stage_6_0_t800;
reg [6-1:0] FSM_fft_64_stage_6_0_t801;
reg [32-1:0] FSM_fft_64_stage_6_0_t802;
reg [6-1:0] FSM_fft_64_stage_6_0_t803;
reg [32-1:0] FSM_fft_64_stage_6_0_t804;
reg [32-1:0] FSM_fft_64_stage_6_0_t805;
reg [6-1:0] FSM_fft_64_stage_6_0_t806;
reg [32-1:0] FSM_fft_64_stage_6_0_t807;
reg [33-1:0] FSM_fft_64_stage_6_0_t808;
reg [32-1:0] FSM_fft_64_stage_6_0_t809;
reg [2048-1:0] FSM_fft_64_stage_6_0_t810;
reg [32-1:0] FSM_fft_64_stage_6_0_t811;
reg [6-1:0] FSM_fft_64_stage_6_0_t812;
reg [32-1:0] FSM_fft_64_stage_6_0_t813;
reg [6-1:0] FSM_fft_64_stage_6_0_t814;
reg [32-1:0] FSM_fft_64_stage_6_0_t815;
reg [32-1:0] FSM_fft_64_stage_6_0_t816;
reg [6-1:0] FSM_fft_64_stage_6_0_t817;
reg [32-1:0] FSM_fft_64_stage_6_0_t818;
reg [2048-1:0] FSM_fft_64_stage_6_0_t819;
reg [32-1:0] FSM_fft_64_stage_6_0_t820;
reg [6-1:0] FSM_fft_64_stage_6_0_t821;
reg [32-1:0] FSM_fft_64_stage_6_0_t822;
reg [6-1:0] FSM_fft_64_stage_6_0_t823;
reg [32-1:0] FSM_fft_64_stage_6_0_t824;
reg [32-1:0] FSM_fft_64_stage_6_0_t825;
reg [6-1:0] FSM_fft_64_stage_6_0_t826;
reg [32-1:0] FSM_fft_64_stage_6_0_t827;
reg [33-1:0] FSM_fft_64_stage_6_0_t828;
reg [32-1:0] FSM_fft_64_stage_6_0_t829;
reg [2048-1:0] FSM_fft_64_stage_6_0_t830;
reg [32-1:0] FSM_fft_64_stage_6_0_t831;
reg [6-1:0] FSM_fft_64_stage_6_0_t832;
reg [32-1:0] FSM_fft_64_stage_6_0_t833;
reg [6-1:0] FSM_fft_64_stage_6_0_t834;
reg [32-1:0] FSM_fft_64_stage_6_0_t835;
reg [32-1:0] FSM_fft_64_stage_6_0_t836;
reg [6-1:0] FSM_fft_64_stage_6_0_t837;
reg [32-1:0] FSM_fft_64_stage_6_0_t838;
reg [2048-1:0] FSM_fft_64_stage_6_0_t839;
reg [32-1:0] FSM_fft_64_stage_6_0_t840;
reg [6-1:0] FSM_fft_64_stage_6_0_t841;
reg [32-1:0] FSM_fft_64_stage_6_0_t842;
reg [6-1:0] FSM_fft_64_stage_6_0_t843;
reg [32-1:0] FSM_fft_64_stage_6_0_t844;
reg [32-1:0] FSM_fft_64_stage_6_0_t845;
reg [6-1:0] FSM_fft_64_stage_6_0_t846;
reg [32-1:0] FSM_fft_64_stage_6_0_t847;
reg [33-1:0] FSM_fft_64_stage_6_0_t848;
reg [32-1:0] FSM_fft_64_stage_6_0_t849;
reg [2048-1:0] FSM_fft_64_stage_6_0_t850;
reg [32-1:0] FSM_fft_64_stage_6_0_t851;
reg [6-1:0] FSM_fft_64_stage_6_0_t852;
reg [32-1:0] FSM_fft_64_stage_6_0_t853;
reg [6-1:0] FSM_fft_64_stage_6_0_t854;
reg [32-1:0] FSM_fft_64_stage_6_0_t855;
reg [32-1:0] FSM_fft_64_stage_6_0_t856;
reg [6-1:0] FSM_fft_64_stage_6_0_t857;
reg [32-1:0] FSM_fft_64_stage_6_0_t858;
reg [2048-1:0] FSM_fft_64_stage_6_0_t859;
reg [32-1:0] FSM_fft_64_stage_6_0_t860;
reg [6-1:0] FSM_fft_64_stage_6_0_t861;
reg [32-1:0] FSM_fft_64_stage_6_0_t862;
reg [6-1:0] FSM_fft_64_stage_6_0_t863;
reg [32-1:0] FSM_fft_64_stage_6_0_t864;
reg [32-1:0] FSM_fft_64_stage_6_0_t865;
reg [6-1:0] FSM_fft_64_stage_6_0_t866;
reg [32-1:0] FSM_fft_64_stage_6_0_t867;
reg [33-1:0] FSM_fft_64_stage_6_0_t868;
reg [32-1:0] FSM_fft_64_stage_6_0_t869;
reg [2048-1:0] FSM_fft_64_stage_6_0_t870;
reg [32-1:0] FSM_fft_64_stage_6_0_t871;
reg [6-1:0] FSM_fft_64_stage_6_0_t872;
reg [32-1:0] FSM_fft_64_stage_6_0_t873;
reg [6-1:0] FSM_fft_64_stage_6_0_t874;
reg [32-1:0] FSM_fft_64_stage_6_0_t875;
reg [32-1:0] FSM_fft_64_stage_6_0_t876;
reg [6-1:0] FSM_fft_64_stage_6_0_t877;
reg [32-1:0] FSM_fft_64_stage_6_0_t878;
reg [2048-1:0] FSM_fft_64_stage_6_0_t879;
reg [32-1:0] FSM_fft_64_stage_6_0_t880;
reg [6-1:0] FSM_fft_64_stage_6_0_t881;
reg [32-1:0] FSM_fft_64_stage_6_0_t882;
reg [6-1:0] FSM_fft_64_stage_6_0_t883;
reg [32-1:0] FSM_fft_64_stage_6_0_t884;
reg [32-1:0] FSM_fft_64_stage_6_0_t885;
reg [6-1:0] FSM_fft_64_stage_6_0_t886;
reg [32-1:0] FSM_fft_64_stage_6_0_t887;
reg [33-1:0] FSM_fft_64_stage_6_0_t888;
reg [32-1:0] FSM_fft_64_stage_6_0_t889;
reg [2048-1:0] FSM_fft_64_stage_6_0_t890;
reg [32-1:0] FSM_fft_64_stage_6_0_t891;
reg [6-1:0] FSM_fft_64_stage_6_0_t892;
reg [32-1:0] FSM_fft_64_stage_6_0_t893;
reg [6-1:0] FSM_fft_64_stage_6_0_t894;
reg [32-1:0] FSM_fft_64_stage_6_0_t895;
reg [32-1:0] FSM_fft_64_stage_6_0_t896;
reg [6-1:0] FSM_fft_64_stage_6_0_t897;
reg [32-1:0] FSM_fft_64_stage_6_0_t898;
reg [2048-1:0] FSM_fft_64_stage_6_0_t899;
reg [32-1:0] FSM_fft_64_stage_6_0_t900;
reg [6-1:0] FSM_fft_64_stage_6_0_t901;
reg [32-1:0] FSM_fft_64_stage_6_0_t902;
reg [6-1:0] FSM_fft_64_stage_6_0_t903;
reg [32-1:0] FSM_fft_64_stage_6_0_t904;
reg [32-1:0] FSM_fft_64_stage_6_0_t905;
reg [6-1:0] FSM_fft_64_stage_6_0_t906;
reg [32-1:0] FSM_fft_64_stage_6_0_t907;
reg [33-1:0] FSM_fft_64_stage_6_0_t908;
reg [32-1:0] FSM_fft_64_stage_6_0_t909;
reg [2048-1:0] FSM_fft_64_stage_6_0_t910;
reg [32-1:0] FSM_fft_64_stage_6_0_t911;
reg [6-1:0] FSM_fft_64_stage_6_0_t912;
reg [32-1:0] FSM_fft_64_stage_6_0_t913;
reg [6-1:0] FSM_fft_64_stage_6_0_t914;
reg [32-1:0] FSM_fft_64_stage_6_0_t915;
reg [32-1:0] FSM_fft_64_stage_6_0_t916;
reg [6-1:0] FSM_fft_64_stage_6_0_t917;
reg [32-1:0] FSM_fft_64_stage_6_0_t918;
reg [2048-1:0] FSM_fft_64_stage_6_0_t919;
reg [32-1:0] FSM_fft_64_stage_6_0_t920;
reg [6-1:0] FSM_fft_64_stage_6_0_t921;
reg [32-1:0] FSM_fft_64_stage_6_0_t922;
reg [6-1:0] FSM_fft_64_stage_6_0_t923;
reg [32-1:0] FSM_fft_64_stage_6_0_t924;
reg [32-1:0] FSM_fft_64_stage_6_0_t925;
reg [6-1:0] FSM_fft_64_stage_6_0_t926;
reg [32-1:0] FSM_fft_64_stage_6_0_t927;
reg [33-1:0] FSM_fft_64_stage_6_0_t928;
reg [32-1:0] FSM_fft_64_stage_6_0_t929;
reg [2048-1:0] FSM_fft_64_stage_6_0_t930;
reg [32-1:0] FSM_fft_64_stage_6_0_t931;
reg [6-1:0] FSM_fft_64_stage_6_0_t932;
reg [32-1:0] FSM_fft_64_stage_6_0_t933;
reg [6-1:0] FSM_fft_64_stage_6_0_t934;
reg [32-1:0] FSM_fft_64_stage_6_0_t935;
reg [32-1:0] FSM_fft_64_stage_6_0_t936;
reg [6-1:0] FSM_fft_64_stage_6_0_t937;
reg [32-1:0] FSM_fft_64_stage_6_0_t938;
reg [2048-1:0] FSM_fft_64_stage_6_0_t939;
reg [32-1:0] FSM_fft_64_stage_6_0_t940;
reg [6-1:0] FSM_fft_64_stage_6_0_t941;
reg [32-1:0] FSM_fft_64_stage_6_0_t942;
reg [6-1:0] FSM_fft_64_stage_6_0_t943;
reg [32-1:0] FSM_fft_64_stage_6_0_t944;
reg [32-1:0] FSM_fft_64_stage_6_0_t945;
reg [6-1:0] FSM_fft_64_stage_6_0_t946;
reg [32-1:0] FSM_fft_64_stage_6_0_t947;
reg [33-1:0] FSM_fft_64_stage_6_0_t948;
reg [32-1:0] FSM_fft_64_stage_6_0_t949;
reg [2048-1:0] FSM_fft_64_stage_6_0_t950;
reg [32-1:0] FSM_fft_64_stage_6_0_t951;
reg [6-1:0] FSM_fft_64_stage_6_0_t952;
reg [32-1:0] FSM_fft_64_stage_6_0_t953;
reg [6-1:0] FSM_fft_64_stage_6_0_t954;
reg [32-1:0] FSM_fft_64_stage_6_0_t955;
reg [32-1:0] FSM_fft_64_stage_6_0_t956;
reg [6-1:0] FSM_fft_64_stage_6_0_t957;
reg [32-1:0] FSM_fft_64_stage_6_0_t958;
reg [2048-1:0] FSM_fft_64_stage_6_0_t959;
reg [32-1:0] FSM_fft_64_stage_6_0_t960;
reg [6-1:0] FSM_fft_64_stage_6_0_t961;
reg [32-1:0] FSM_fft_64_stage_6_0_t962;
reg [6-1:0] FSM_fft_64_stage_6_0_t963;
reg [32-1:0] FSM_fft_64_stage_6_0_t964;
reg [32-1:0] FSM_fft_64_stage_6_0_t965;
reg [6-1:0] FSM_fft_64_stage_6_0_t966;
reg [32-1:0] FSM_fft_64_stage_6_0_t967;
reg [33-1:0] FSM_fft_64_stage_6_0_t968;
reg [32-1:0] FSM_fft_64_stage_6_0_t969;
reg [2048-1:0] FSM_fft_64_stage_6_0_t970;
reg [32-1:0] FSM_fft_64_stage_6_0_t971;
reg [6-1:0] FSM_fft_64_stage_6_0_t972;
reg [32-1:0] FSM_fft_64_stage_6_0_t973;
reg [6-1:0] FSM_fft_64_stage_6_0_t974;
reg [32-1:0] FSM_fft_64_stage_6_0_t975;
reg [32-1:0] FSM_fft_64_stage_6_0_t976;
reg [6-1:0] FSM_fft_64_stage_6_0_t977;
reg [32-1:0] FSM_fft_64_stage_6_0_t978;
reg [2048-1:0] FSM_fft_64_stage_6_0_t979;
reg [32-1:0] FSM_fft_64_stage_6_0_t980;
reg [6-1:0] FSM_fft_64_stage_6_0_t981;
reg [32-1:0] FSM_fft_64_stage_6_0_t982;
reg [6-1:0] FSM_fft_64_stage_6_0_t983;
reg [32-1:0] FSM_fft_64_stage_6_0_t984;
reg [32-1:0] FSM_fft_64_stage_6_0_t985;
reg [6-1:0] FSM_fft_64_stage_6_0_t986;
reg [32-1:0] FSM_fft_64_stage_6_0_t987;
reg [33-1:0] FSM_fft_64_stage_6_0_t988;
reg [32-1:0] FSM_fft_64_stage_6_0_t989;
reg [2048-1:0] FSM_fft_64_stage_6_0_t990;
reg [32-1:0] FSM_fft_64_stage_6_0_t991;
reg [6-1:0] FSM_fft_64_stage_6_0_t992;
reg [32-1:0] FSM_fft_64_stage_6_0_t993;
reg [6-1:0] FSM_fft_64_stage_6_0_t994;
reg [32-1:0] FSM_fft_64_stage_6_0_t995;
reg [32-1:0] FSM_fft_64_stage_6_0_t996;
reg [6-1:0] FSM_fft_64_stage_6_0_t997;
reg [32-1:0] FSM_fft_64_stage_6_0_t998;
reg [2048-1:0] FSM_fft_64_stage_6_0_t999;
reg [32-1:0] FSM_fft_64_stage_6_0_t1000;
reg [6-1:0] FSM_fft_64_stage_6_0_t1001;
reg [32-1:0] FSM_fft_64_stage_6_0_t1002;
reg [6-1:0] FSM_fft_64_stage_6_0_t1003;
reg [32-1:0] FSM_fft_64_stage_6_0_t1004;
reg [32-1:0] FSM_fft_64_stage_6_0_t1005;
reg [6-1:0] FSM_fft_64_stage_6_0_t1006;
reg [32-1:0] FSM_fft_64_stage_6_0_t1007;
reg [33-1:0] FSM_fft_64_stage_6_0_t1008;
reg [32-1:0] FSM_fft_64_stage_6_0_t1009;
reg [2048-1:0] FSM_fft_64_stage_6_0_t1010;
reg [32-1:0] FSM_fft_64_stage_6_0_t1011;
reg [6-1:0] FSM_fft_64_stage_6_0_t1012;
reg [32-1:0] FSM_fft_64_stage_6_0_t1013;
reg [6-1:0] FSM_fft_64_stage_6_0_t1014;
reg [32-1:0] FSM_fft_64_stage_6_0_t1015;
reg [32-1:0] FSM_fft_64_stage_6_0_t1016;
reg [6-1:0] FSM_fft_64_stage_6_0_t1017;
reg [32-1:0] FSM_fft_64_stage_6_0_t1018;
reg [2048-1:0] FSM_fft_64_stage_6_0_t1019;
reg [32-1:0] FSM_fft_64_stage_6_0_t1020;
reg [6-1:0] FSM_fft_64_stage_6_0_t1021;
reg [32-1:0] FSM_fft_64_stage_6_0_t1022;
reg [6-1:0] FSM_fft_64_stage_6_0_t1023;
reg [32-1:0] FSM_fft_64_stage_6_0_t1024;
reg [32-1:0] FSM_fft_64_stage_6_0_t1025;
reg [6-1:0] FSM_fft_64_stage_6_0_t1026;
reg [32-1:0] FSM_fft_64_stage_6_0_t1027;
reg [33-1:0] FSM_fft_64_stage_6_0_t1028;
reg [32-1:0] FSM_fft_64_stage_6_0_t1029;
reg [2048-1:0] FSM_fft_64_stage_6_0_t1030;
reg [32-1:0] FSM_fft_64_stage_6_0_t1031;
reg [6-1:0] FSM_fft_64_stage_6_0_t1032;
reg [32-1:0] FSM_fft_64_stage_6_0_t1033;
reg [6-1:0] FSM_fft_64_stage_6_0_t1034;
reg [32-1:0] FSM_fft_64_stage_6_0_t1035;
reg [32-1:0] FSM_fft_64_stage_6_0_t1036;
reg [6-1:0] FSM_fft_64_stage_6_0_t1037;
reg [32-1:0] FSM_fft_64_stage_6_0_t1038;
reg [2048-1:0] FSM_fft_64_stage_6_0_t1039;
reg [32-1:0] FSM_fft_64_stage_6_0_t1040;
reg [6-1:0] FSM_fft_64_stage_6_0_t1041;
reg [32-1:0] FSM_fft_64_stage_6_0_t1042;
reg [6-1:0] FSM_fft_64_stage_6_0_t1043;
reg [32-1:0] FSM_fft_64_stage_6_0_t1044;
reg [32-1:0] FSM_fft_64_stage_6_0_t1045;
reg [6-1:0] FSM_fft_64_stage_6_0_t1046;
reg [32-1:0] FSM_fft_64_stage_6_0_t1047;
reg [33-1:0] FSM_fft_64_stage_6_0_t1048;
reg [32-1:0] FSM_fft_64_stage_6_0_t1049;
reg [2048-1:0] FSM_fft_64_stage_6_0_t1050;
reg [32-1:0] FSM_fft_64_stage_6_0_t1051;
reg [6-1:0] FSM_fft_64_stage_6_0_t1052;
reg [32-1:0] FSM_fft_64_stage_6_0_t1053;
reg [6-1:0] FSM_fft_64_stage_6_0_t1054;
reg [32-1:0] FSM_fft_64_stage_6_0_t1055;
reg [32-1:0] FSM_fft_64_stage_6_0_t1056;
reg [6-1:0] FSM_fft_64_stage_6_0_t1057;
reg [32-1:0] FSM_fft_64_stage_6_0_t1058;
reg [2048-1:0] FSM_fft_64_stage_6_0_t1059;
reg [32-1:0] FSM_fft_64_stage_6_0_t1060;
reg [6-1:0] FSM_fft_64_stage_6_0_t1061;
reg [32-1:0] FSM_fft_64_stage_6_0_t1062;
reg [6-1:0] FSM_fft_64_stage_6_0_t1063;
reg [32-1:0] FSM_fft_64_stage_6_0_t1064;
reg [32-1:0] FSM_fft_64_stage_6_0_t1065;
reg [6-1:0] FSM_fft_64_stage_6_0_t1066;
reg [32-1:0] FSM_fft_64_stage_6_0_t1067;
reg [33-1:0] FSM_fft_64_stage_6_0_t1068;
reg [32-1:0] FSM_fft_64_stage_6_0_t1069;
reg [2048-1:0] FSM_fft_64_stage_6_0_t1070;
reg [32-1:0] FSM_fft_64_stage_6_0_t1071;
reg [6-1:0] FSM_fft_64_stage_6_0_t1072;
reg [32-1:0] FSM_fft_64_stage_6_0_t1073;
reg [6-1:0] FSM_fft_64_stage_6_0_t1074;
reg [32-1:0] FSM_fft_64_stage_6_0_t1075;
reg [32-1:0] FSM_fft_64_stage_6_0_t1076;
reg [6-1:0] FSM_fft_64_stage_6_0_t1077;
reg [32-1:0] FSM_fft_64_stage_6_0_t1078;
reg [2048-1:0] FSM_fft_64_stage_6_0_t1079;
reg [32-1:0] FSM_fft_64_stage_6_0_t1080;
reg [6-1:0] FSM_fft_64_stage_6_0_t1081;
reg [32-1:0] FSM_fft_64_stage_6_0_t1082;
reg [6-1:0] FSM_fft_64_stage_6_0_t1083;
reg [32-1:0] FSM_fft_64_stage_6_0_t1084;
reg [32-1:0] FSM_fft_64_stage_6_0_t1085;
reg [6-1:0] FSM_fft_64_stage_6_0_t1086;
reg [32-1:0] FSM_fft_64_stage_6_0_t1087;
reg [33-1:0] FSM_fft_64_stage_6_0_t1088;
reg [32-1:0] FSM_fft_64_stage_6_0_t1089;
reg [2048-1:0] FSM_fft_64_stage_6_0_t1090;
reg [32-1:0] FSM_fft_64_stage_6_0_t1091;
reg [6-1:0] FSM_fft_64_stage_6_0_t1092;
reg [32-1:0] FSM_fft_64_stage_6_0_t1093;
reg [6-1:0] FSM_fft_64_stage_6_0_t1094;
reg [32-1:0] FSM_fft_64_stage_6_0_t1095;
reg [32-1:0] FSM_fft_64_stage_6_0_t1096;
reg [6-1:0] FSM_fft_64_stage_6_0_t1097;
reg [32-1:0] FSM_fft_64_stage_6_0_t1098;
reg [2048-1:0] FSM_fft_64_stage_6_0_t1099;
reg [32-1:0] FSM_fft_64_stage_6_0_t1100;
reg [6-1:0] FSM_fft_64_stage_6_0_t1101;
reg [32-1:0] FSM_fft_64_stage_6_0_t1102;
reg [6-1:0] FSM_fft_64_stage_6_0_t1103;
reg [32-1:0] FSM_fft_64_stage_6_0_t1104;
reg [32-1:0] FSM_fft_64_stage_6_0_t1105;
reg [6-1:0] FSM_fft_64_stage_6_0_t1106;
reg [32-1:0] FSM_fft_64_stage_6_0_t1107;
reg [33-1:0] FSM_fft_64_stage_6_0_t1108;
reg [32-1:0] FSM_fft_64_stage_6_0_t1109;
reg [2048-1:0] FSM_fft_64_stage_6_0_t1110;
reg [32-1:0] FSM_fft_64_stage_6_0_t1111;
reg [6-1:0] FSM_fft_64_stage_6_0_t1112;
reg [32-1:0] FSM_fft_64_stage_6_0_t1113;
reg [6-1:0] FSM_fft_64_stage_6_0_t1114;
reg [32-1:0] FSM_fft_64_stage_6_0_t1115;
reg [32-1:0] FSM_fft_64_stage_6_0_t1116;
reg [6-1:0] FSM_fft_64_stage_6_0_t1117;
reg [32-1:0] FSM_fft_64_stage_6_0_t1118;
reg [2048-1:0] FSM_fft_64_stage_6_0_t1119;
reg [32-1:0] FSM_fft_64_stage_6_0_t1120;
reg [6-1:0] FSM_fft_64_stage_6_0_t1121;
reg [32-1:0] FSM_fft_64_stage_6_0_t1122;
reg [6-1:0] FSM_fft_64_stage_6_0_t1123;
reg [32-1:0] FSM_fft_64_stage_6_0_t1124;
reg [32-1:0] FSM_fft_64_stage_6_0_t1125;
reg [6-1:0] FSM_fft_64_stage_6_0_t1126;
reg [32-1:0] FSM_fft_64_stage_6_0_t1127;
reg [33-1:0] FSM_fft_64_stage_6_0_t1128;
reg [32-1:0] FSM_fft_64_stage_6_0_t1129;
reg [2048-1:0] FSM_fft_64_stage_6_0_t1130;
reg [32-1:0] FSM_fft_64_stage_6_0_t1131;
reg [6-1:0] FSM_fft_64_stage_6_0_t1132;
reg [32-1:0] FSM_fft_64_stage_6_0_t1133;
reg [6-1:0] FSM_fft_64_stage_6_0_t1134;
reg [32-1:0] FSM_fft_64_stage_6_0_t1135;
reg [32-1:0] FSM_fft_64_stage_6_0_t1136;
reg [6-1:0] FSM_fft_64_stage_6_0_t1137;
reg [32-1:0] FSM_fft_64_stage_6_0_t1138;
reg [2048-1:0] FSM_fft_64_stage_6_0_t1139;
reg [32-1:0] FSM_fft_64_stage_6_0_t1140;
reg [6-1:0] FSM_fft_64_stage_6_0_t1141;
reg [32-1:0] FSM_fft_64_stage_6_0_t1142;
reg [6-1:0] FSM_fft_64_stage_6_0_t1143;
reg [32-1:0] FSM_fft_64_stage_6_0_t1144;
reg [32-1:0] FSM_fft_64_stage_6_0_t1145;
reg [6-1:0] FSM_fft_64_stage_6_0_t1146;
reg [32-1:0] FSM_fft_64_stage_6_0_t1147;
reg [33-1:0] FSM_fft_64_stage_6_0_t1148;
reg [32-1:0] FSM_fft_64_stage_6_0_t1149;
reg [2048-1:0] FSM_fft_64_stage_6_0_t1150;
reg [32-1:0] FSM_fft_64_stage_6_0_t1151;
reg [6-1:0] FSM_fft_64_stage_6_0_t1152;
reg [32-1:0] FSM_fft_64_stage_6_0_t1153;
reg [6-1:0] FSM_fft_64_stage_6_0_t1154;
reg [32-1:0] FSM_fft_64_stage_6_0_t1155;
reg [32-1:0] FSM_fft_64_stage_6_0_t1156;
reg [6-1:0] FSM_fft_64_stage_6_0_t1157;
reg [32-1:0] FSM_fft_64_stage_6_0_t1158;
reg [2048-1:0] FSM_fft_64_stage_6_0_t1159;
reg [32-1:0] FSM_fft_64_stage_6_0_t1160;
reg [6-1:0] FSM_fft_64_stage_6_0_t1161;
reg [32-1:0] FSM_fft_64_stage_6_0_t1162;
reg [6-1:0] FSM_fft_64_stage_6_0_t1163;
reg [32-1:0] FSM_fft_64_stage_6_0_t1164;
reg [32-1:0] FSM_fft_64_stage_6_0_t1165;
reg [6-1:0] FSM_fft_64_stage_6_0_t1166;
reg [32-1:0] FSM_fft_64_stage_6_0_t1167;
reg [33-1:0] FSM_fft_64_stage_6_0_t1168;
reg [32-1:0] FSM_fft_64_stage_6_0_t1169;
reg [2048-1:0] FSM_fft_64_stage_6_0_t1170;
reg [32-1:0] FSM_fft_64_stage_6_0_t1171;
reg [6-1:0] FSM_fft_64_stage_6_0_t1172;
reg [32-1:0] FSM_fft_64_stage_6_0_t1173;
reg [6-1:0] FSM_fft_64_stage_6_0_t1174;
reg [32-1:0] FSM_fft_64_stage_6_0_t1175;
reg [32-1:0] FSM_fft_64_stage_6_0_t1176;
reg [6-1:0] FSM_fft_64_stage_6_0_t1177;
reg [32-1:0] FSM_fft_64_stage_6_0_t1178;
reg [2048-1:0] FSM_fft_64_stage_6_0_t1179;
reg [32-1:0] FSM_fft_64_stage_6_0_t1180;
reg [6-1:0] FSM_fft_64_stage_6_0_t1181;
reg [32-1:0] FSM_fft_64_stage_6_0_t1182;
reg [6-1:0] FSM_fft_64_stage_6_0_t1183;
reg [32-1:0] FSM_fft_64_stage_6_0_t1184;
reg [32-1:0] FSM_fft_64_stage_6_0_t1185;
reg [6-1:0] FSM_fft_64_stage_6_0_t1186;
reg [32-1:0] FSM_fft_64_stage_6_0_t1187;
reg [33-1:0] FSM_fft_64_stage_6_0_t1188;
reg [32-1:0] FSM_fft_64_stage_6_0_t1189;
reg [2048-1:0] FSM_fft_64_stage_6_0_t1190;
reg [32-1:0] FSM_fft_64_stage_6_0_t1191;
reg [6-1:0] FSM_fft_64_stage_6_0_t1192;
reg [32-1:0] FSM_fft_64_stage_6_0_t1193;
reg [6-1:0] FSM_fft_64_stage_6_0_t1194;
reg [32-1:0] FSM_fft_64_stage_6_0_t1195;
reg [32-1:0] FSM_fft_64_stage_6_0_t1196;
reg [6-1:0] FSM_fft_64_stage_6_0_t1197;
reg [32-1:0] FSM_fft_64_stage_6_0_t1198;
reg [2048-1:0] FSM_fft_64_stage_6_0_t1199;
reg [32-1:0] FSM_fft_64_stage_6_0_t1200;
reg [6-1:0] FSM_fft_64_stage_6_0_t1201;
reg [32-1:0] FSM_fft_64_stage_6_0_t1202;
reg [6-1:0] FSM_fft_64_stage_6_0_t1203;
reg [32-1:0] FSM_fft_64_stage_6_0_t1204;
reg [32-1:0] FSM_fft_64_stage_6_0_t1205;
reg [6-1:0] FSM_fft_64_stage_6_0_t1206;
reg [32-1:0] FSM_fft_64_stage_6_0_t1207;
reg [33-1:0] FSM_fft_64_stage_6_0_t1208;
reg [32-1:0] FSM_fft_64_stage_6_0_t1209;
reg [2048-1:0] FSM_fft_64_stage_6_0_t1210;
reg [32-1:0] FSM_fft_64_stage_6_0_t1211;
reg [6-1:0] FSM_fft_64_stage_6_0_t1212;
reg [32-1:0] FSM_fft_64_stage_6_0_t1213;
reg [6-1:0] FSM_fft_64_stage_6_0_t1214;
reg [32-1:0] FSM_fft_64_stage_6_0_t1215;
reg [32-1:0] FSM_fft_64_stage_6_0_t1216;
reg [6-1:0] FSM_fft_64_stage_6_0_t1217;
reg [32-1:0] FSM_fft_64_stage_6_0_t1218;
reg [2048-1:0] FSM_fft_64_stage_6_0_t1219;
reg [32-1:0] FSM_fft_64_stage_6_0_t1220;
reg [6-1:0] FSM_fft_64_stage_6_0_t1221;
reg [32-1:0] FSM_fft_64_stage_6_0_t1222;
reg [6-1:0] FSM_fft_64_stage_6_0_t1223;
reg [32-1:0] FSM_fft_64_stage_6_0_t1224;
reg [32-1:0] FSM_fft_64_stage_6_0_t1225;
reg [6-1:0] FSM_fft_64_stage_6_0_t1226;
reg [32-1:0] FSM_fft_64_stage_6_0_t1227;
reg [33-1:0] FSM_fft_64_stage_6_0_t1228;
reg [32-1:0] FSM_fft_64_stage_6_0_t1229;
reg [2048-1:0] FSM_fft_64_stage_6_0_t1230;
reg [32-1:0] FSM_fft_64_stage_6_0_t1231;
reg [6-1:0] FSM_fft_64_stage_6_0_t1232;
reg [32-1:0] FSM_fft_64_stage_6_0_t1233;
reg [6-1:0] FSM_fft_64_stage_6_0_t1234;
reg [32-1:0] FSM_fft_64_stage_6_0_t1235;
reg [32-1:0] FSM_fft_64_stage_6_0_t1236;
reg [6-1:0] FSM_fft_64_stage_6_0_t1237;
reg [32-1:0] FSM_fft_64_stage_6_0_t1238;
reg [2048-1:0] FSM_fft_64_stage_6_0_t1239;
reg [32-1:0] FSM_fft_64_stage_6_0_t1240;
reg [6-1:0] FSM_fft_64_stage_6_0_t1241;
reg [32-1:0] FSM_fft_64_stage_6_0_t1242;
reg [6-1:0] FSM_fft_64_stage_6_0_t1243;
reg [32-1:0] FSM_fft_64_stage_6_0_t1244;
reg [32-1:0] FSM_fft_64_stage_6_0_t1245;
reg [6-1:0] FSM_fft_64_stage_6_0_t1246;
reg [32-1:0] FSM_fft_64_stage_6_0_t1247;
reg [33-1:0] FSM_fft_64_stage_6_0_t1248;
reg [32-1:0] FSM_fft_64_stage_6_0_t1249;
reg [2048-1:0] FSM_fft_64_stage_6_0_t1250;
reg [32-1:0] FSM_fft_64_stage_6_0_t1251;
reg [6-1:0] FSM_fft_64_stage_6_0_t1252;
reg [32-1:0] FSM_fft_64_stage_6_0_t1253;
reg [6-1:0] FSM_fft_64_stage_6_0_t1254;
reg [32-1:0] FSM_fft_64_stage_6_0_t1255;
reg [32-1:0] FSM_fft_64_stage_6_0_t1256;
reg [6-1:0] FSM_fft_64_stage_6_0_t1257;
reg [32-1:0] FSM_fft_64_stage_6_0_t1258;
reg [2048-1:0] FSM_fft_64_stage_6_0_t1259;
reg [32-1:0] FSM_fft_64_stage_6_0_t1260;
reg [6-1:0] FSM_fft_64_stage_6_0_t1261;
reg [32-1:0] FSM_fft_64_stage_6_0_t1262;
reg [6-1:0] FSM_fft_64_stage_6_0_t1263;
reg [32-1:0] FSM_fft_64_stage_6_0_t1264;
reg [32-1:0] FSM_fft_64_stage_6_0_t1265;
reg [6-1:0] FSM_fft_64_stage_6_0_t1266;
reg [32-1:0] FSM_fft_64_stage_6_0_t1267;
reg [33-1:0] FSM_fft_64_stage_6_0_t1268;
reg [32-1:0] FSM_fft_64_stage_6_0_t1269;
reg [2048-1:0] FSM_fft_64_stage_6_0_t1270;
reg [32-1:0] FSM_fft_64_stage_6_0_t1271;
reg [6-1:0] FSM_fft_64_stage_6_0_t1272;
reg [32-1:0] FSM_fft_64_stage_6_0_t1273;
reg [6-1:0] FSM_fft_64_stage_6_0_t1274;
reg [32-1:0] FSM_fft_64_stage_6_0_t1275;
reg [32-1:0] FSM_fft_64_stage_6_0_t1276;
reg [6-1:0] FSM_fft_64_stage_6_0_t1277;
reg [32-1:0] FSM_fft_64_stage_6_0_t1278;
reg [2048-1:0] FSM_fft_64_stage_6_0_t1279;

assign FSM_fft_64_stage_6_0_out_valid = 1'b1;
/*
    Wiring by fft_64_stage_6
*/
assign i_ready = FSM_fft_64_stage_6_0_in_ready;
assign o_data_out_real = FSM_fft_64_stage_6_0_t639;
assign o_data_out_imag = FSM_fft_64_stage_6_0_t1279;
assign o_valid = FSM_fft_64_stage_6_0_out_valid;
/* End wiring by fft_64_stage_6 */

initial begin
    FSM_fft_64_stage_6_0_t0 = 32'b0;
    FSM_fft_64_stage_6_0_t1 = FSM_fft_64_stage_6_0_t0[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t2 = 32'b0;
    FSM_fft_64_stage_6_0_t3 = FSM_fft_64_stage_6_0_t2[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t4 = i_data_in_real[FSM_fft_64_stage_6_0_t3 * 32 +: 32];
    FSM_fft_64_stage_6_0_t5 = 32'b00000000000000000000000000100000;
    FSM_fft_64_stage_6_0_t6 = FSM_fft_64_stage_6_0_t5[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t7 = i_data_in_real[FSM_fft_64_stage_6_0_t6 * 32 +: 32];
    FSM_fft_64_stage_6_0_t8 = FSM_fft_64_stage_6_0_t4 + FSM_fft_64_stage_6_0_t7;
    FSM_fft_64_stage_6_0_t9 = FSM_fft_64_stage_6_0_t8[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t10 = i_data_in_real;
    FSM_fft_64_stage_6_0_t10[FSM_fft_64_stage_6_0_t1 * 32 +: 32] = FSM_fft_64_stage_6_0_t9;
    FSM_fft_64_stage_6_0_t11 = 32'b00000000000000000000000000100000;
    FSM_fft_64_stage_6_0_t12 = FSM_fft_64_stage_6_0_t11[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t13 = 32'b0;
    FSM_fft_64_stage_6_0_t14 = FSM_fft_64_stage_6_0_t13[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t15 = i_data_in_real[FSM_fft_64_stage_6_0_t14 * 32 +: 32];
    FSM_fft_64_stage_6_0_t16 = 32'b00000000000000000000000000100000;
    FSM_fft_64_stage_6_0_t17 = FSM_fft_64_stage_6_0_t16[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t18 = i_data_in_real[FSM_fft_64_stage_6_0_t17 * 32 +: 32];
    FSM_fft_64_stage_6_0_t19 = FSM_fft_64_stage_6_0_t10;
    FSM_fft_64_stage_6_0_t19[FSM_fft_64_stage_6_0_t12 * 32 +: 32] = FSM_fft_64_stage_6_0_t15 - FSM_fft_64_stage_6_0_t18;
    FSM_fft_64_stage_6_0_t20 = 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_6_0_t21 = FSM_fft_64_stage_6_0_t20[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t22 = 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_6_0_t23 = FSM_fft_64_stage_6_0_t22[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t24 = i_data_in_real[FSM_fft_64_stage_6_0_t23 * 32 +: 32];
    FSM_fft_64_stage_6_0_t25 = 32'b00000000000000000000000000100001;
    FSM_fft_64_stage_6_0_t26 = FSM_fft_64_stage_6_0_t25[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t27 = i_data_in_real[FSM_fft_64_stage_6_0_t26 * 32 +: 32];
    FSM_fft_64_stage_6_0_t28 = FSM_fft_64_stage_6_0_t24 + FSM_fft_64_stage_6_0_t27;
    FSM_fft_64_stage_6_0_t29 = FSM_fft_64_stage_6_0_t28[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t30 = FSM_fft_64_stage_6_0_t19;
    FSM_fft_64_stage_6_0_t30[FSM_fft_64_stage_6_0_t21 * 32 +: 32] = FSM_fft_64_stage_6_0_t29;
    FSM_fft_64_stage_6_0_t31 = 32'b00000000000000000000000000100001;
    FSM_fft_64_stage_6_0_t32 = FSM_fft_64_stage_6_0_t31[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t33 = 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_6_0_t34 = FSM_fft_64_stage_6_0_t33[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t35 = i_data_in_real[FSM_fft_64_stage_6_0_t34 * 32 +: 32];
    FSM_fft_64_stage_6_0_t36 = 32'b00000000000000000000000000100001;
    FSM_fft_64_stage_6_0_t37 = FSM_fft_64_stage_6_0_t36[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t38 = i_data_in_real[FSM_fft_64_stage_6_0_t37 * 32 +: 32];
    FSM_fft_64_stage_6_0_t39 = FSM_fft_64_stage_6_0_t30;
    FSM_fft_64_stage_6_0_t39[FSM_fft_64_stage_6_0_t32 * 32 +: 32] = FSM_fft_64_stage_6_0_t35 - FSM_fft_64_stage_6_0_t38;
    FSM_fft_64_stage_6_0_t40 = 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_6_0_t41 = FSM_fft_64_stage_6_0_t40[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t42 = 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_6_0_t43 = FSM_fft_64_stage_6_0_t42[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t44 = i_data_in_real[FSM_fft_64_stage_6_0_t43 * 32 +: 32];
    FSM_fft_64_stage_6_0_t45 = 32'b00000000000000000000000000100010;
    FSM_fft_64_stage_6_0_t46 = FSM_fft_64_stage_6_0_t45[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t47 = i_data_in_real[FSM_fft_64_stage_6_0_t46 * 32 +: 32];
    FSM_fft_64_stage_6_0_t48 = FSM_fft_64_stage_6_0_t44 + FSM_fft_64_stage_6_0_t47;
    FSM_fft_64_stage_6_0_t49 = FSM_fft_64_stage_6_0_t48[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t50 = FSM_fft_64_stage_6_0_t39;
    FSM_fft_64_stage_6_0_t50[FSM_fft_64_stage_6_0_t41 * 32 +: 32] = FSM_fft_64_stage_6_0_t49;
    FSM_fft_64_stage_6_0_t51 = 32'b00000000000000000000000000100010;
    FSM_fft_64_stage_6_0_t52 = FSM_fft_64_stage_6_0_t51[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t53 = 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_6_0_t54 = FSM_fft_64_stage_6_0_t53[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t55 = i_data_in_real[FSM_fft_64_stage_6_0_t54 * 32 +: 32];
    FSM_fft_64_stage_6_0_t56 = 32'b00000000000000000000000000100010;
    FSM_fft_64_stage_6_0_t57 = FSM_fft_64_stage_6_0_t56[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t58 = i_data_in_real[FSM_fft_64_stage_6_0_t57 * 32 +: 32];
    FSM_fft_64_stage_6_0_t59 = FSM_fft_64_stage_6_0_t50;
    FSM_fft_64_stage_6_0_t59[FSM_fft_64_stage_6_0_t52 * 32 +: 32] = FSM_fft_64_stage_6_0_t55 - FSM_fft_64_stage_6_0_t58;
    FSM_fft_64_stage_6_0_t60 = 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_6_0_t61 = FSM_fft_64_stage_6_0_t60[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t62 = 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_6_0_t63 = FSM_fft_64_stage_6_0_t62[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t64 = i_data_in_real[FSM_fft_64_stage_6_0_t63 * 32 +: 32];
    FSM_fft_64_stage_6_0_t65 = 32'b00000000000000000000000000100011;
    FSM_fft_64_stage_6_0_t66 = FSM_fft_64_stage_6_0_t65[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t67 = i_data_in_real[FSM_fft_64_stage_6_0_t66 * 32 +: 32];
    FSM_fft_64_stage_6_0_t68 = FSM_fft_64_stage_6_0_t64 + FSM_fft_64_stage_6_0_t67;
    FSM_fft_64_stage_6_0_t69 = FSM_fft_64_stage_6_0_t68[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t70 = FSM_fft_64_stage_6_0_t59;
    FSM_fft_64_stage_6_0_t70[FSM_fft_64_stage_6_0_t61 * 32 +: 32] = FSM_fft_64_stage_6_0_t69;
    FSM_fft_64_stage_6_0_t71 = 32'b00000000000000000000000000100011;
    FSM_fft_64_stage_6_0_t72 = FSM_fft_64_stage_6_0_t71[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t73 = 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_6_0_t74 = FSM_fft_64_stage_6_0_t73[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t75 = i_data_in_real[FSM_fft_64_stage_6_0_t74 * 32 +: 32];
    FSM_fft_64_stage_6_0_t76 = 32'b00000000000000000000000000100011;
    FSM_fft_64_stage_6_0_t77 = FSM_fft_64_stage_6_0_t76[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t78 = i_data_in_real[FSM_fft_64_stage_6_0_t77 * 32 +: 32];
    FSM_fft_64_stage_6_0_t79 = FSM_fft_64_stage_6_0_t70;
    FSM_fft_64_stage_6_0_t79[FSM_fft_64_stage_6_0_t72 * 32 +: 32] = FSM_fft_64_stage_6_0_t75 - FSM_fft_64_stage_6_0_t78;
    FSM_fft_64_stage_6_0_t80 = 32'b00000000000000000000000000000100;
    FSM_fft_64_stage_6_0_t81 = FSM_fft_64_stage_6_0_t80[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t82 = 32'b00000000000000000000000000000100;
    FSM_fft_64_stage_6_0_t83 = FSM_fft_64_stage_6_0_t82[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t84 = i_data_in_real[FSM_fft_64_stage_6_0_t83 * 32 +: 32];
    FSM_fft_64_stage_6_0_t85 = 32'b00000000000000000000000000100100;
    FSM_fft_64_stage_6_0_t86 = FSM_fft_64_stage_6_0_t85[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t87 = i_data_in_real[FSM_fft_64_stage_6_0_t86 * 32 +: 32];
    FSM_fft_64_stage_6_0_t88 = FSM_fft_64_stage_6_0_t84 + FSM_fft_64_stage_6_0_t87;
    FSM_fft_64_stage_6_0_t89 = FSM_fft_64_stage_6_0_t88[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t90 = FSM_fft_64_stage_6_0_t79;
    FSM_fft_64_stage_6_0_t90[FSM_fft_64_stage_6_0_t81 * 32 +: 32] = FSM_fft_64_stage_6_0_t89;
    FSM_fft_64_stage_6_0_t91 = 32'b00000000000000000000000000100100;
    FSM_fft_64_stage_6_0_t92 = FSM_fft_64_stage_6_0_t91[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t93 = 32'b00000000000000000000000000000100;
    FSM_fft_64_stage_6_0_t94 = FSM_fft_64_stage_6_0_t93[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t95 = i_data_in_real[FSM_fft_64_stage_6_0_t94 * 32 +: 32];
    FSM_fft_64_stage_6_0_t96 = 32'b00000000000000000000000000100100;
    FSM_fft_64_stage_6_0_t97 = FSM_fft_64_stage_6_0_t96[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t98 = i_data_in_real[FSM_fft_64_stage_6_0_t97 * 32 +: 32];
    FSM_fft_64_stage_6_0_t99 = FSM_fft_64_stage_6_0_t90;
    FSM_fft_64_stage_6_0_t99[FSM_fft_64_stage_6_0_t92 * 32 +: 32] = FSM_fft_64_stage_6_0_t95 - FSM_fft_64_stage_6_0_t98;
    FSM_fft_64_stage_6_0_t100 = 32'b00000000000000000000000000000101;
    FSM_fft_64_stage_6_0_t101 = FSM_fft_64_stage_6_0_t100[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t102 = 32'b00000000000000000000000000000101;
    FSM_fft_64_stage_6_0_t103 = FSM_fft_64_stage_6_0_t102[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t104 = i_data_in_real[FSM_fft_64_stage_6_0_t103 * 32 +: 32];
    FSM_fft_64_stage_6_0_t105 = 32'b00000000000000000000000000100101;
    FSM_fft_64_stage_6_0_t106 = FSM_fft_64_stage_6_0_t105[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t107 = i_data_in_real[FSM_fft_64_stage_6_0_t106 * 32 +: 32];
    FSM_fft_64_stage_6_0_t108 = FSM_fft_64_stage_6_0_t104 + FSM_fft_64_stage_6_0_t107;
    FSM_fft_64_stage_6_0_t109 = FSM_fft_64_stage_6_0_t108[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t110 = FSM_fft_64_stage_6_0_t99;
    FSM_fft_64_stage_6_0_t110[FSM_fft_64_stage_6_0_t101 * 32 +: 32] = FSM_fft_64_stage_6_0_t109;
    FSM_fft_64_stage_6_0_t111 = 32'b00000000000000000000000000100101;
    FSM_fft_64_stage_6_0_t112 = FSM_fft_64_stage_6_0_t111[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t113 = 32'b00000000000000000000000000000101;
    FSM_fft_64_stage_6_0_t114 = FSM_fft_64_stage_6_0_t113[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t115 = i_data_in_real[FSM_fft_64_stage_6_0_t114 * 32 +: 32];
    FSM_fft_64_stage_6_0_t116 = 32'b00000000000000000000000000100101;
    FSM_fft_64_stage_6_0_t117 = FSM_fft_64_stage_6_0_t116[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t118 = i_data_in_real[FSM_fft_64_stage_6_0_t117 * 32 +: 32];
    FSM_fft_64_stage_6_0_t119 = FSM_fft_64_stage_6_0_t110;
    FSM_fft_64_stage_6_0_t119[FSM_fft_64_stage_6_0_t112 * 32 +: 32] = FSM_fft_64_stage_6_0_t115 - FSM_fft_64_stage_6_0_t118;
    FSM_fft_64_stage_6_0_t120 = 32'b00000000000000000000000000000110;
    FSM_fft_64_stage_6_0_t121 = FSM_fft_64_stage_6_0_t120[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t122 = 32'b00000000000000000000000000000110;
    FSM_fft_64_stage_6_0_t123 = FSM_fft_64_stage_6_0_t122[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t124 = i_data_in_real[FSM_fft_64_stage_6_0_t123 * 32 +: 32];
    FSM_fft_64_stage_6_0_t125 = 32'b00000000000000000000000000100110;
    FSM_fft_64_stage_6_0_t126 = FSM_fft_64_stage_6_0_t125[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t127 = i_data_in_real[FSM_fft_64_stage_6_0_t126 * 32 +: 32];
    FSM_fft_64_stage_6_0_t128 = FSM_fft_64_stage_6_0_t124 + FSM_fft_64_stage_6_0_t127;
    FSM_fft_64_stage_6_0_t129 = FSM_fft_64_stage_6_0_t128[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t130 = FSM_fft_64_stage_6_0_t119;
    FSM_fft_64_stage_6_0_t130[FSM_fft_64_stage_6_0_t121 * 32 +: 32] = FSM_fft_64_stage_6_0_t129;
    FSM_fft_64_stage_6_0_t131 = 32'b00000000000000000000000000100110;
    FSM_fft_64_stage_6_0_t132 = FSM_fft_64_stage_6_0_t131[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t133 = 32'b00000000000000000000000000000110;
    FSM_fft_64_stage_6_0_t134 = FSM_fft_64_stage_6_0_t133[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t135 = i_data_in_real[FSM_fft_64_stage_6_0_t134 * 32 +: 32];
    FSM_fft_64_stage_6_0_t136 = 32'b00000000000000000000000000100110;
    FSM_fft_64_stage_6_0_t137 = FSM_fft_64_stage_6_0_t136[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t138 = i_data_in_real[FSM_fft_64_stage_6_0_t137 * 32 +: 32];
    FSM_fft_64_stage_6_0_t139 = FSM_fft_64_stage_6_0_t130;
    FSM_fft_64_stage_6_0_t139[FSM_fft_64_stage_6_0_t132 * 32 +: 32] = FSM_fft_64_stage_6_0_t135 - FSM_fft_64_stage_6_0_t138;
    FSM_fft_64_stage_6_0_t140 = 32'b00000000000000000000000000000111;
    FSM_fft_64_stage_6_0_t141 = FSM_fft_64_stage_6_0_t140[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t142 = 32'b00000000000000000000000000000111;
    FSM_fft_64_stage_6_0_t143 = FSM_fft_64_stage_6_0_t142[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t144 = i_data_in_real[FSM_fft_64_stage_6_0_t143 * 32 +: 32];
    FSM_fft_64_stage_6_0_t145 = 32'b00000000000000000000000000100111;
    FSM_fft_64_stage_6_0_t146 = FSM_fft_64_stage_6_0_t145[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t147 = i_data_in_real[FSM_fft_64_stage_6_0_t146 * 32 +: 32];
    FSM_fft_64_stage_6_0_t148 = FSM_fft_64_stage_6_0_t144 + FSM_fft_64_stage_6_0_t147;
    FSM_fft_64_stage_6_0_t149 = FSM_fft_64_stage_6_0_t148[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t150 = FSM_fft_64_stage_6_0_t139;
    FSM_fft_64_stage_6_0_t150[FSM_fft_64_stage_6_0_t141 * 32 +: 32] = FSM_fft_64_stage_6_0_t149;
    FSM_fft_64_stage_6_0_t151 = 32'b00000000000000000000000000100111;
    FSM_fft_64_stage_6_0_t152 = FSM_fft_64_stage_6_0_t151[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t153 = 32'b00000000000000000000000000000111;
    FSM_fft_64_stage_6_0_t154 = FSM_fft_64_stage_6_0_t153[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t155 = i_data_in_real[FSM_fft_64_stage_6_0_t154 * 32 +: 32];
    FSM_fft_64_stage_6_0_t156 = 32'b00000000000000000000000000100111;
    FSM_fft_64_stage_6_0_t157 = FSM_fft_64_stage_6_0_t156[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t158 = i_data_in_real[FSM_fft_64_stage_6_0_t157 * 32 +: 32];
    FSM_fft_64_stage_6_0_t159 = FSM_fft_64_stage_6_0_t150;
    FSM_fft_64_stage_6_0_t159[FSM_fft_64_stage_6_0_t152 * 32 +: 32] = FSM_fft_64_stage_6_0_t155 - FSM_fft_64_stage_6_0_t158;
    FSM_fft_64_stage_6_0_t160 = 32'b00000000000000000000000000001000;
    FSM_fft_64_stage_6_0_t161 = FSM_fft_64_stage_6_0_t160[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t162 = 32'b00000000000000000000000000001000;
    FSM_fft_64_stage_6_0_t163 = FSM_fft_64_stage_6_0_t162[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t164 = i_data_in_real[FSM_fft_64_stage_6_0_t163 * 32 +: 32];
    FSM_fft_64_stage_6_0_t165 = 32'b00000000000000000000000000101000;
    FSM_fft_64_stage_6_0_t166 = FSM_fft_64_stage_6_0_t165[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t167 = i_data_in_real[FSM_fft_64_stage_6_0_t166 * 32 +: 32];
    FSM_fft_64_stage_6_0_t168 = FSM_fft_64_stage_6_0_t164 + FSM_fft_64_stage_6_0_t167;
    FSM_fft_64_stage_6_0_t169 = FSM_fft_64_stage_6_0_t168[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t170 = FSM_fft_64_stage_6_0_t159;
    FSM_fft_64_stage_6_0_t170[FSM_fft_64_stage_6_0_t161 * 32 +: 32] = FSM_fft_64_stage_6_0_t169;
    FSM_fft_64_stage_6_0_t171 = 32'b00000000000000000000000000101000;
    FSM_fft_64_stage_6_0_t172 = FSM_fft_64_stage_6_0_t171[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t173 = 32'b00000000000000000000000000001000;
    FSM_fft_64_stage_6_0_t174 = FSM_fft_64_stage_6_0_t173[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t175 = i_data_in_real[FSM_fft_64_stage_6_0_t174 * 32 +: 32];
    FSM_fft_64_stage_6_0_t176 = 32'b00000000000000000000000000101000;
    FSM_fft_64_stage_6_0_t177 = FSM_fft_64_stage_6_0_t176[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t178 = i_data_in_real[FSM_fft_64_stage_6_0_t177 * 32 +: 32];
    FSM_fft_64_stage_6_0_t179 = FSM_fft_64_stage_6_0_t170;
    FSM_fft_64_stage_6_0_t179[FSM_fft_64_stage_6_0_t172 * 32 +: 32] = FSM_fft_64_stage_6_0_t175 - FSM_fft_64_stage_6_0_t178;
    FSM_fft_64_stage_6_0_t180 = 32'b00000000000000000000000000001001;
    FSM_fft_64_stage_6_0_t181 = FSM_fft_64_stage_6_0_t180[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t182 = 32'b00000000000000000000000000001001;
    FSM_fft_64_stage_6_0_t183 = FSM_fft_64_stage_6_0_t182[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t184 = i_data_in_real[FSM_fft_64_stage_6_0_t183 * 32 +: 32];
    FSM_fft_64_stage_6_0_t185 = 32'b00000000000000000000000000101001;
    FSM_fft_64_stage_6_0_t186 = FSM_fft_64_stage_6_0_t185[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t187 = i_data_in_real[FSM_fft_64_stage_6_0_t186 * 32 +: 32];
    FSM_fft_64_stage_6_0_t188 = FSM_fft_64_stage_6_0_t184 + FSM_fft_64_stage_6_0_t187;
    FSM_fft_64_stage_6_0_t189 = FSM_fft_64_stage_6_0_t188[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t190 = FSM_fft_64_stage_6_0_t179;
    FSM_fft_64_stage_6_0_t190[FSM_fft_64_stage_6_0_t181 * 32 +: 32] = FSM_fft_64_stage_6_0_t189;
    FSM_fft_64_stage_6_0_t191 = 32'b00000000000000000000000000101001;
    FSM_fft_64_stage_6_0_t192 = FSM_fft_64_stage_6_0_t191[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t193 = 32'b00000000000000000000000000001001;
    FSM_fft_64_stage_6_0_t194 = FSM_fft_64_stage_6_0_t193[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t195 = i_data_in_real[FSM_fft_64_stage_6_0_t194 * 32 +: 32];
    FSM_fft_64_stage_6_0_t196 = 32'b00000000000000000000000000101001;
    FSM_fft_64_stage_6_0_t197 = FSM_fft_64_stage_6_0_t196[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t198 = i_data_in_real[FSM_fft_64_stage_6_0_t197 * 32 +: 32];
    FSM_fft_64_stage_6_0_t199 = FSM_fft_64_stage_6_0_t190;
    FSM_fft_64_stage_6_0_t199[FSM_fft_64_stage_6_0_t192 * 32 +: 32] = FSM_fft_64_stage_6_0_t195 - FSM_fft_64_stage_6_0_t198;
    FSM_fft_64_stage_6_0_t200 = 32'b00000000000000000000000000001010;
    FSM_fft_64_stage_6_0_t201 = FSM_fft_64_stage_6_0_t200[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t202 = 32'b00000000000000000000000000001010;
    FSM_fft_64_stage_6_0_t203 = FSM_fft_64_stage_6_0_t202[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t204 = i_data_in_real[FSM_fft_64_stage_6_0_t203 * 32 +: 32];
    FSM_fft_64_stage_6_0_t205 = 32'b00000000000000000000000000101010;
    FSM_fft_64_stage_6_0_t206 = FSM_fft_64_stage_6_0_t205[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t207 = i_data_in_real[FSM_fft_64_stage_6_0_t206 * 32 +: 32];
    FSM_fft_64_stage_6_0_t208 = FSM_fft_64_stage_6_0_t204 + FSM_fft_64_stage_6_0_t207;
    FSM_fft_64_stage_6_0_t209 = FSM_fft_64_stage_6_0_t208[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t210 = FSM_fft_64_stage_6_0_t199;
    FSM_fft_64_stage_6_0_t210[FSM_fft_64_stage_6_0_t201 * 32 +: 32] = FSM_fft_64_stage_6_0_t209;
    FSM_fft_64_stage_6_0_t211 = 32'b00000000000000000000000000101010;
    FSM_fft_64_stage_6_0_t212 = FSM_fft_64_stage_6_0_t211[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t213 = 32'b00000000000000000000000000001010;
    FSM_fft_64_stage_6_0_t214 = FSM_fft_64_stage_6_0_t213[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t215 = i_data_in_real[FSM_fft_64_stage_6_0_t214 * 32 +: 32];
    FSM_fft_64_stage_6_0_t216 = 32'b00000000000000000000000000101010;
    FSM_fft_64_stage_6_0_t217 = FSM_fft_64_stage_6_0_t216[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t218 = i_data_in_real[FSM_fft_64_stage_6_0_t217 * 32 +: 32];
    FSM_fft_64_stage_6_0_t219 = FSM_fft_64_stage_6_0_t210;
    FSM_fft_64_stage_6_0_t219[FSM_fft_64_stage_6_0_t212 * 32 +: 32] = FSM_fft_64_stage_6_0_t215 - FSM_fft_64_stage_6_0_t218;
    FSM_fft_64_stage_6_0_t220 = 32'b00000000000000000000000000001011;
    FSM_fft_64_stage_6_0_t221 = FSM_fft_64_stage_6_0_t220[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t222 = 32'b00000000000000000000000000001011;
    FSM_fft_64_stage_6_0_t223 = FSM_fft_64_stage_6_0_t222[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t224 = i_data_in_real[FSM_fft_64_stage_6_0_t223 * 32 +: 32];
    FSM_fft_64_stage_6_0_t225 = 32'b00000000000000000000000000101011;
    FSM_fft_64_stage_6_0_t226 = FSM_fft_64_stage_6_0_t225[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t227 = i_data_in_real[FSM_fft_64_stage_6_0_t226 * 32 +: 32];
    FSM_fft_64_stage_6_0_t228 = FSM_fft_64_stage_6_0_t224 + FSM_fft_64_stage_6_0_t227;
    FSM_fft_64_stage_6_0_t229 = FSM_fft_64_stage_6_0_t228[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t230 = FSM_fft_64_stage_6_0_t219;
    FSM_fft_64_stage_6_0_t230[FSM_fft_64_stage_6_0_t221 * 32 +: 32] = FSM_fft_64_stage_6_0_t229;
    FSM_fft_64_stage_6_0_t231 = 32'b00000000000000000000000000101011;
    FSM_fft_64_stage_6_0_t232 = FSM_fft_64_stage_6_0_t231[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t233 = 32'b00000000000000000000000000001011;
    FSM_fft_64_stage_6_0_t234 = FSM_fft_64_stage_6_0_t233[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t235 = i_data_in_real[FSM_fft_64_stage_6_0_t234 * 32 +: 32];
    FSM_fft_64_stage_6_0_t236 = 32'b00000000000000000000000000101011;
    FSM_fft_64_stage_6_0_t237 = FSM_fft_64_stage_6_0_t236[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t238 = i_data_in_real[FSM_fft_64_stage_6_0_t237 * 32 +: 32];
    FSM_fft_64_stage_6_0_t239 = FSM_fft_64_stage_6_0_t230;
    FSM_fft_64_stage_6_0_t239[FSM_fft_64_stage_6_0_t232 * 32 +: 32] = FSM_fft_64_stage_6_0_t235 - FSM_fft_64_stage_6_0_t238;
    FSM_fft_64_stage_6_0_t240 = 32'b00000000000000000000000000001100;
    FSM_fft_64_stage_6_0_t241 = FSM_fft_64_stage_6_0_t240[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t242 = 32'b00000000000000000000000000001100;
    FSM_fft_64_stage_6_0_t243 = FSM_fft_64_stage_6_0_t242[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t244 = i_data_in_real[FSM_fft_64_stage_6_0_t243 * 32 +: 32];
    FSM_fft_64_stage_6_0_t245 = 32'b00000000000000000000000000101100;
    FSM_fft_64_stage_6_0_t246 = FSM_fft_64_stage_6_0_t245[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t247 = i_data_in_real[FSM_fft_64_stage_6_0_t246 * 32 +: 32];
    FSM_fft_64_stage_6_0_t248 = FSM_fft_64_stage_6_0_t244 + FSM_fft_64_stage_6_0_t247;
    FSM_fft_64_stage_6_0_t249 = FSM_fft_64_stage_6_0_t248[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t250 = FSM_fft_64_stage_6_0_t239;
    FSM_fft_64_stage_6_0_t250[FSM_fft_64_stage_6_0_t241 * 32 +: 32] = FSM_fft_64_stage_6_0_t249;
    FSM_fft_64_stage_6_0_t251 = 32'b00000000000000000000000000101100;
    FSM_fft_64_stage_6_0_t252 = FSM_fft_64_stage_6_0_t251[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t253 = 32'b00000000000000000000000000001100;
    FSM_fft_64_stage_6_0_t254 = FSM_fft_64_stage_6_0_t253[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t255 = i_data_in_real[FSM_fft_64_stage_6_0_t254 * 32 +: 32];
    FSM_fft_64_stage_6_0_t256 = 32'b00000000000000000000000000101100;
    FSM_fft_64_stage_6_0_t257 = FSM_fft_64_stage_6_0_t256[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t258 = i_data_in_real[FSM_fft_64_stage_6_0_t257 * 32 +: 32];
    FSM_fft_64_stage_6_0_t259 = FSM_fft_64_stage_6_0_t250;
    FSM_fft_64_stage_6_0_t259[FSM_fft_64_stage_6_0_t252 * 32 +: 32] = FSM_fft_64_stage_6_0_t255 - FSM_fft_64_stage_6_0_t258;
    FSM_fft_64_stage_6_0_t260 = 32'b00000000000000000000000000001101;
    FSM_fft_64_stage_6_0_t261 = FSM_fft_64_stage_6_0_t260[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t262 = 32'b00000000000000000000000000001101;
    FSM_fft_64_stage_6_0_t263 = FSM_fft_64_stage_6_0_t262[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t264 = i_data_in_real[FSM_fft_64_stage_6_0_t263 * 32 +: 32];
    FSM_fft_64_stage_6_0_t265 = 32'b00000000000000000000000000101101;
    FSM_fft_64_stage_6_0_t266 = FSM_fft_64_stage_6_0_t265[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t267 = i_data_in_real[FSM_fft_64_stage_6_0_t266 * 32 +: 32];
    FSM_fft_64_stage_6_0_t268 = FSM_fft_64_stage_6_0_t264 + FSM_fft_64_stage_6_0_t267;
    FSM_fft_64_stage_6_0_t269 = FSM_fft_64_stage_6_0_t268[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t270 = FSM_fft_64_stage_6_0_t259;
    FSM_fft_64_stage_6_0_t270[FSM_fft_64_stage_6_0_t261 * 32 +: 32] = FSM_fft_64_stage_6_0_t269;
    FSM_fft_64_stage_6_0_t271 = 32'b00000000000000000000000000101101;
    FSM_fft_64_stage_6_0_t272 = FSM_fft_64_stage_6_0_t271[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t273 = 32'b00000000000000000000000000001101;
    FSM_fft_64_stage_6_0_t274 = FSM_fft_64_stage_6_0_t273[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t275 = i_data_in_real[FSM_fft_64_stage_6_0_t274 * 32 +: 32];
    FSM_fft_64_stage_6_0_t276 = 32'b00000000000000000000000000101101;
    FSM_fft_64_stage_6_0_t277 = FSM_fft_64_stage_6_0_t276[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t278 = i_data_in_real[FSM_fft_64_stage_6_0_t277 * 32 +: 32];
    FSM_fft_64_stage_6_0_t279 = FSM_fft_64_stage_6_0_t270;
    FSM_fft_64_stage_6_0_t279[FSM_fft_64_stage_6_0_t272 * 32 +: 32] = FSM_fft_64_stage_6_0_t275 - FSM_fft_64_stage_6_0_t278;
    FSM_fft_64_stage_6_0_t280 = 32'b00000000000000000000000000001110;
    FSM_fft_64_stage_6_0_t281 = FSM_fft_64_stage_6_0_t280[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t282 = 32'b00000000000000000000000000001110;
    FSM_fft_64_stage_6_0_t283 = FSM_fft_64_stage_6_0_t282[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t284 = i_data_in_real[FSM_fft_64_stage_6_0_t283 * 32 +: 32];
    FSM_fft_64_stage_6_0_t285 = 32'b00000000000000000000000000101110;
    FSM_fft_64_stage_6_0_t286 = FSM_fft_64_stage_6_0_t285[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t287 = i_data_in_real[FSM_fft_64_stage_6_0_t286 * 32 +: 32];
    FSM_fft_64_stage_6_0_t288 = FSM_fft_64_stage_6_0_t284 + FSM_fft_64_stage_6_0_t287;
    FSM_fft_64_stage_6_0_t289 = FSM_fft_64_stage_6_0_t288[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t290 = FSM_fft_64_stage_6_0_t279;
    FSM_fft_64_stage_6_0_t290[FSM_fft_64_stage_6_0_t281 * 32 +: 32] = FSM_fft_64_stage_6_0_t289;
    FSM_fft_64_stage_6_0_t291 = 32'b00000000000000000000000000101110;
    FSM_fft_64_stage_6_0_t292 = FSM_fft_64_stage_6_0_t291[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t293 = 32'b00000000000000000000000000001110;
    FSM_fft_64_stage_6_0_t294 = FSM_fft_64_stage_6_0_t293[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t295 = i_data_in_real[FSM_fft_64_stage_6_0_t294 * 32 +: 32];
    FSM_fft_64_stage_6_0_t296 = 32'b00000000000000000000000000101110;
    FSM_fft_64_stage_6_0_t297 = FSM_fft_64_stage_6_0_t296[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t298 = i_data_in_real[FSM_fft_64_stage_6_0_t297 * 32 +: 32];
    FSM_fft_64_stage_6_0_t299 = FSM_fft_64_stage_6_0_t290;
    FSM_fft_64_stage_6_0_t299[FSM_fft_64_stage_6_0_t292 * 32 +: 32] = FSM_fft_64_stage_6_0_t295 - FSM_fft_64_stage_6_0_t298;
    FSM_fft_64_stage_6_0_t300 = 32'b00000000000000000000000000001111;
    FSM_fft_64_stage_6_0_t301 = FSM_fft_64_stage_6_0_t300[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t302 = 32'b00000000000000000000000000001111;
    FSM_fft_64_stage_6_0_t303 = FSM_fft_64_stage_6_0_t302[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t304 = i_data_in_real[FSM_fft_64_stage_6_0_t303 * 32 +: 32];
    FSM_fft_64_stage_6_0_t305 = 32'b00000000000000000000000000101111;
    FSM_fft_64_stage_6_0_t306 = FSM_fft_64_stage_6_0_t305[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t307 = i_data_in_real[FSM_fft_64_stage_6_0_t306 * 32 +: 32];
    FSM_fft_64_stage_6_0_t308 = FSM_fft_64_stage_6_0_t304 + FSM_fft_64_stage_6_0_t307;
    FSM_fft_64_stage_6_0_t309 = FSM_fft_64_stage_6_0_t308[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t310 = FSM_fft_64_stage_6_0_t299;
    FSM_fft_64_stage_6_0_t310[FSM_fft_64_stage_6_0_t301 * 32 +: 32] = FSM_fft_64_stage_6_0_t309;
    FSM_fft_64_stage_6_0_t311 = 32'b00000000000000000000000000101111;
    FSM_fft_64_stage_6_0_t312 = FSM_fft_64_stage_6_0_t311[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t313 = 32'b00000000000000000000000000001111;
    FSM_fft_64_stage_6_0_t314 = FSM_fft_64_stage_6_0_t313[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t315 = i_data_in_real[FSM_fft_64_stage_6_0_t314 * 32 +: 32];
    FSM_fft_64_stage_6_0_t316 = 32'b00000000000000000000000000101111;
    FSM_fft_64_stage_6_0_t317 = FSM_fft_64_stage_6_0_t316[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t318 = i_data_in_real[FSM_fft_64_stage_6_0_t317 * 32 +: 32];
    FSM_fft_64_stage_6_0_t319 = FSM_fft_64_stage_6_0_t310;
    FSM_fft_64_stage_6_0_t319[FSM_fft_64_stage_6_0_t312 * 32 +: 32] = FSM_fft_64_stage_6_0_t315 - FSM_fft_64_stage_6_0_t318;
    FSM_fft_64_stage_6_0_t320 = 32'b00000000000000000000000000010000;
    FSM_fft_64_stage_6_0_t321 = FSM_fft_64_stage_6_0_t320[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t322 = 32'b00000000000000000000000000010000;
    FSM_fft_64_stage_6_0_t323 = FSM_fft_64_stage_6_0_t322[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t324 = i_data_in_real[FSM_fft_64_stage_6_0_t323 * 32 +: 32];
    FSM_fft_64_stage_6_0_t325 = 32'b00000000000000000000000000110000;
    FSM_fft_64_stage_6_0_t326 = FSM_fft_64_stage_6_0_t325[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t327 = i_data_in_real[FSM_fft_64_stage_6_0_t326 * 32 +: 32];
    FSM_fft_64_stage_6_0_t328 = FSM_fft_64_stage_6_0_t324 + FSM_fft_64_stage_6_0_t327;
    FSM_fft_64_stage_6_0_t329 = FSM_fft_64_stage_6_0_t328[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t330 = FSM_fft_64_stage_6_0_t319;
    FSM_fft_64_stage_6_0_t330[FSM_fft_64_stage_6_0_t321 * 32 +: 32] = FSM_fft_64_stage_6_0_t329;
    FSM_fft_64_stage_6_0_t331 = 32'b00000000000000000000000000110000;
    FSM_fft_64_stage_6_0_t332 = FSM_fft_64_stage_6_0_t331[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t333 = 32'b00000000000000000000000000010000;
    FSM_fft_64_stage_6_0_t334 = FSM_fft_64_stage_6_0_t333[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t335 = i_data_in_real[FSM_fft_64_stage_6_0_t334 * 32 +: 32];
    FSM_fft_64_stage_6_0_t336 = 32'b00000000000000000000000000110000;
    FSM_fft_64_stage_6_0_t337 = FSM_fft_64_stage_6_0_t336[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t338 = i_data_in_real[FSM_fft_64_stage_6_0_t337 * 32 +: 32];
    FSM_fft_64_stage_6_0_t339 = FSM_fft_64_stage_6_0_t330;
    FSM_fft_64_stage_6_0_t339[FSM_fft_64_stage_6_0_t332 * 32 +: 32] = FSM_fft_64_stage_6_0_t335 - FSM_fft_64_stage_6_0_t338;
    FSM_fft_64_stage_6_0_t340 = 32'b00000000000000000000000000010001;
    FSM_fft_64_stage_6_0_t341 = FSM_fft_64_stage_6_0_t340[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t342 = 32'b00000000000000000000000000010001;
    FSM_fft_64_stage_6_0_t343 = FSM_fft_64_stage_6_0_t342[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t344 = i_data_in_real[FSM_fft_64_stage_6_0_t343 * 32 +: 32];
    FSM_fft_64_stage_6_0_t345 = 32'b00000000000000000000000000110001;
    FSM_fft_64_stage_6_0_t346 = FSM_fft_64_stage_6_0_t345[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t347 = i_data_in_real[FSM_fft_64_stage_6_0_t346 * 32 +: 32];
    FSM_fft_64_stage_6_0_t348 = FSM_fft_64_stage_6_0_t344 + FSM_fft_64_stage_6_0_t347;
    FSM_fft_64_stage_6_0_t349 = FSM_fft_64_stage_6_0_t348[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t350 = FSM_fft_64_stage_6_0_t339;
    FSM_fft_64_stage_6_0_t350[FSM_fft_64_stage_6_0_t341 * 32 +: 32] = FSM_fft_64_stage_6_0_t349;
    FSM_fft_64_stage_6_0_t351 = 32'b00000000000000000000000000110001;
    FSM_fft_64_stage_6_0_t352 = FSM_fft_64_stage_6_0_t351[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t353 = 32'b00000000000000000000000000010001;
    FSM_fft_64_stage_6_0_t354 = FSM_fft_64_stage_6_0_t353[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t355 = i_data_in_real[FSM_fft_64_stage_6_0_t354 * 32 +: 32];
    FSM_fft_64_stage_6_0_t356 = 32'b00000000000000000000000000110001;
    FSM_fft_64_stage_6_0_t357 = FSM_fft_64_stage_6_0_t356[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t358 = i_data_in_real[FSM_fft_64_stage_6_0_t357 * 32 +: 32];
    FSM_fft_64_stage_6_0_t359 = FSM_fft_64_stage_6_0_t350;
    FSM_fft_64_stage_6_0_t359[FSM_fft_64_stage_6_0_t352 * 32 +: 32] = FSM_fft_64_stage_6_0_t355 - FSM_fft_64_stage_6_0_t358;
    FSM_fft_64_stage_6_0_t360 = 32'b00000000000000000000000000010010;
    FSM_fft_64_stage_6_0_t361 = FSM_fft_64_stage_6_0_t360[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t362 = 32'b00000000000000000000000000010010;
    FSM_fft_64_stage_6_0_t363 = FSM_fft_64_stage_6_0_t362[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t364 = i_data_in_real[FSM_fft_64_stage_6_0_t363 * 32 +: 32];
    FSM_fft_64_stage_6_0_t365 = 32'b00000000000000000000000000110010;
    FSM_fft_64_stage_6_0_t366 = FSM_fft_64_stage_6_0_t365[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t367 = i_data_in_real[FSM_fft_64_stage_6_0_t366 * 32 +: 32];
    FSM_fft_64_stage_6_0_t368 = FSM_fft_64_stage_6_0_t364 + FSM_fft_64_stage_6_0_t367;
    FSM_fft_64_stage_6_0_t369 = FSM_fft_64_stage_6_0_t368[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t370 = FSM_fft_64_stage_6_0_t359;
    FSM_fft_64_stage_6_0_t370[FSM_fft_64_stage_6_0_t361 * 32 +: 32] = FSM_fft_64_stage_6_0_t369;
    FSM_fft_64_stage_6_0_t371 = 32'b00000000000000000000000000110010;
    FSM_fft_64_stage_6_0_t372 = FSM_fft_64_stage_6_0_t371[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t373 = 32'b00000000000000000000000000010010;
    FSM_fft_64_stage_6_0_t374 = FSM_fft_64_stage_6_0_t373[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t375 = i_data_in_real[FSM_fft_64_stage_6_0_t374 * 32 +: 32];
    FSM_fft_64_stage_6_0_t376 = 32'b00000000000000000000000000110010;
    FSM_fft_64_stage_6_0_t377 = FSM_fft_64_stage_6_0_t376[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t378 = i_data_in_real[FSM_fft_64_stage_6_0_t377 * 32 +: 32];
    FSM_fft_64_stage_6_0_t379 = FSM_fft_64_stage_6_0_t370;
    FSM_fft_64_stage_6_0_t379[FSM_fft_64_stage_6_0_t372 * 32 +: 32] = FSM_fft_64_stage_6_0_t375 - FSM_fft_64_stage_6_0_t378;
    FSM_fft_64_stage_6_0_t380 = 32'b00000000000000000000000000010011;
    FSM_fft_64_stage_6_0_t381 = FSM_fft_64_stage_6_0_t380[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t382 = 32'b00000000000000000000000000010011;
    FSM_fft_64_stage_6_0_t383 = FSM_fft_64_stage_6_0_t382[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t384 = i_data_in_real[FSM_fft_64_stage_6_0_t383 * 32 +: 32];
    FSM_fft_64_stage_6_0_t385 = 32'b00000000000000000000000000110011;
    FSM_fft_64_stage_6_0_t386 = FSM_fft_64_stage_6_0_t385[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t387 = i_data_in_real[FSM_fft_64_stage_6_0_t386 * 32 +: 32];
    FSM_fft_64_stage_6_0_t388 = FSM_fft_64_stage_6_0_t384 + FSM_fft_64_stage_6_0_t387;
    FSM_fft_64_stage_6_0_t389 = FSM_fft_64_stage_6_0_t388[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t390 = FSM_fft_64_stage_6_0_t379;
    FSM_fft_64_stage_6_0_t390[FSM_fft_64_stage_6_0_t381 * 32 +: 32] = FSM_fft_64_stage_6_0_t389;
    FSM_fft_64_stage_6_0_t391 = 32'b00000000000000000000000000110011;
    FSM_fft_64_stage_6_0_t392 = FSM_fft_64_stage_6_0_t391[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t393 = 32'b00000000000000000000000000010011;
    FSM_fft_64_stage_6_0_t394 = FSM_fft_64_stage_6_0_t393[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t395 = i_data_in_real[FSM_fft_64_stage_6_0_t394 * 32 +: 32];
    FSM_fft_64_stage_6_0_t396 = 32'b00000000000000000000000000110011;
    FSM_fft_64_stage_6_0_t397 = FSM_fft_64_stage_6_0_t396[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t398 = i_data_in_real[FSM_fft_64_stage_6_0_t397 * 32 +: 32];
    FSM_fft_64_stage_6_0_t399 = FSM_fft_64_stage_6_0_t390;
    FSM_fft_64_stage_6_0_t399[FSM_fft_64_stage_6_0_t392 * 32 +: 32] = FSM_fft_64_stage_6_0_t395 - FSM_fft_64_stage_6_0_t398;
    FSM_fft_64_stage_6_0_t400 = 32'b00000000000000000000000000010100;
    FSM_fft_64_stage_6_0_t401 = FSM_fft_64_stage_6_0_t400[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t402 = 32'b00000000000000000000000000010100;
    FSM_fft_64_stage_6_0_t403 = FSM_fft_64_stage_6_0_t402[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t404 = i_data_in_real[FSM_fft_64_stage_6_0_t403 * 32 +: 32];
    FSM_fft_64_stage_6_0_t405 = 32'b00000000000000000000000000110100;
    FSM_fft_64_stage_6_0_t406 = FSM_fft_64_stage_6_0_t405[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t407 = i_data_in_real[FSM_fft_64_stage_6_0_t406 * 32 +: 32];
    FSM_fft_64_stage_6_0_t408 = FSM_fft_64_stage_6_0_t404 + FSM_fft_64_stage_6_0_t407;
    FSM_fft_64_stage_6_0_t409 = FSM_fft_64_stage_6_0_t408[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t410 = FSM_fft_64_stage_6_0_t399;
    FSM_fft_64_stage_6_0_t410[FSM_fft_64_stage_6_0_t401 * 32 +: 32] = FSM_fft_64_stage_6_0_t409;
    FSM_fft_64_stage_6_0_t411 = 32'b00000000000000000000000000110100;
    FSM_fft_64_stage_6_0_t412 = FSM_fft_64_stage_6_0_t411[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t413 = 32'b00000000000000000000000000010100;
    FSM_fft_64_stage_6_0_t414 = FSM_fft_64_stage_6_0_t413[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t415 = i_data_in_real[FSM_fft_64_stage_6_0_t414 * 32 +: 32];
    FSM_fft_64_stage_6_0_t416 = 32'b00000000000000000000000000110100;
    FSM_fft_64_stage_6_0_t417 = FSM_fft_64_stage_6_0_t416[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t418 = i_data_in_real[FSM_fft_64_stage_6_0_t417 * 32 +: 32];
    FSM_fft_64_stage_6_0_t419 = FSM_fft_64_stage_6_0_t410;
    FSM_fft_64_stage_6_0_t419[FSM_fft_64_stage_6_0_t412 * 32 +: 32] = FSM_fft_64_stage_6_0_t415 - FSM_fft_64_stage_6_0_t418;
    FSM_fft_64_stage_6_0_t420 = 32'b00000000000000000000000000010101;
    FSM_fft_64_stage_6_0_t421 = FSM_fft_64_stage_6_0_t420[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t422 = 32'b00000000000000000000000000010101;
    FSM_fft_64_stage_6_0_t423 = FSM_fft_64_stage_6_0_t422[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t424 = i_data_in_real[FSM_fft_64_stage_6_0_t423 * 32 +: 32];
    FSM_fft_64_stage_6_0_t425 = 32'b00000000000000000000000000110101;
    FSM_fft_64_stage_6_0_t426 = FSM_fft_64_stage_6_0_t425[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t427 = i_data_in_real[FSM_fft_64_stage_6_0_t426 * 32 +: 32];
    FSM_fft_64_stage_6_0_t428 = FSM_fft_64_stage_6_0_t424 + FSM_fft_64_stage_6_0_t427;
    FSM_fft_64_stage_6_0_t429 = FSM_fft_64_stage_6_0_t428[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t430 = FSM_fft_64_stage_6_0_t419;
    FSM_fft_64_stage_6_0_t430[FSM_fft_64_stage_6_0_t421 * 32 +: 32] = FSM_fft_64_stage_6_0_t429;
    FSM_fft_64_stage_6_0_t431 = 32'b00000000000000000000000000110101;
    FSM_fft_64_stage_6_0_t432 = FSM_fft_64_stage_6_0_t431[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t433 = 32'b00000000000000000000000000010101;
    FSM_fft_64_stage_6_0_t434 = FSM_fft_64_stage_6_0_t433[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t435 = i_data_in_real[FSM_fft_64_stage_6_0_t434 * 32 +: 32];
    FSM_fft_64_stage_6_0_t436 = 32'b00000000000000000000000000110101;
    FSM_fft_64_stage_6_0_t437 = FSM_fft_64_stage_6_0_t436[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t438 = i_data_in_real[FSM_fft_64_stage_6_0_t437 * 32 +: 32];
    FSM_fft_64_stage_6_0_t439 = FSM_fft_64_stage_6_0_t430;
    FSM_fft_64_stage_6_0_t439[FSM_fft_64_stage_6_0_t432 * 32 +: 32] = FSM_fft_64_stage_6_0_t435 - FSM_fft_64_stage_6_0_t438;
    FSM_fft_64_stage_6_0_t440 = 32'b00000000000000000000000000010110;
    FSM_fft_64_stage_6_0_t441 = FSM_fft_64_stage_6_0_t440[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t442 = 32'b00000000000000000000000000010110;
    FSM_fft_64_stage_6_0_t443 = FSM_fft_64_stage_6_0_t442[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t444 = i_data_in_real[FSM_fft_64_stage_6_0_t443 * 32 +: 32];
    FSM_fft_64_stage_6_0_t445 = 32'b00000000000000000000000000110110;
    FSM_fft_64_stage_6_0_t446 = FSM_fft_64_stage_6_0_t445[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t447 = i_data_in_real[FSM_fft_64_stage_6_0_t446 * 32 +: 32];
    FSM_fft_64_stage_6_0_t448 = FSM_fft_64_stage_6_0_t444 + FSM_fft_64_stage_6_0_t447;
    FSM_fft_64_stage_6_0_t449 = FSM_fft_64_stage_6_0_t448[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t450 = FSM_fft_64_stage_6_0_t439;
    FSM_fft_64_stage_6_0_t450[FSM_fft_64_stage_6_0_t441 * 32 +: 32] = FSM_fft_64_stage_6_0_t449;
    FSM_fft_64_stage_6_0_t451 = 32'b00000000000000000000000000110110;
    FSM_fft_64_stage_6_0_t452 = FSM_fft_64_stage_6_0_t451[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t453 = 32'b00000000000000000000000000010110;
    FSM_fft_64_stage_6_0_t454 = FSM_fft_64_stage_6_0_t453[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t455 = i_data_in_real[FSM_fft_64_stage_6_0_t454 * 32 +: 32];
    FSM_fft_64_stage_6_0_t456 = 32'b00000000000000000000000000110110;
    FSM_fft_64_stage_6_0_t457 = FSM_fft_64_stage_6_0_t456[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t458 = i_data_in_real[FSM_fft_64_stage_6_0_t457 * 32 +: 32];
    FSM_fft_64_stage_6_0_t459 = FSM_fft_64_stage_6_0_t450;
    FSM_fft_64_stage_6_0_t459[FSM_fft_64_stage_6_0_t452 * 32 +: 32] = FSM_fft_64_stage_6_0_t455 - FSM_fft_64_stage_6_0_t458;
    FSM_fft_64_stage_6_0_t460 = 32'b00000000000000000000000000010111;
    FSM_fft_64_stage_6_0_t461 = FSM_fft_64_stage_6_0_t460[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t462 = 32'b00000000000000000000000000010111;
    FSM_fft_64_stage_6_0_t463 = FSM_fft_64_stage_6_0_t462[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t464 = i_data_in_real[FSM_fft_64_stage_6_0_t463 * 32 +: 32];
    FSM_fft_64_stage_6_0_t465 = 32'b00000000000000000000000000110111;
    FSM_fft_64_stage_6_0_t466 = FSM_fft_64_stage_6_0_t465[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t467 = i_data_in_real[FSM_fft_64_stage_6_0_t466 * 32 +: 32];
    FSM_fft_64_stage_6_0_t468 = FSM_fft_64_stage_6_0_t464 + FSM_fft_64_stage_6_0_t467;
    FSM_fft_64_stage_6_0_t469 = FSM_fft_64_stage_6_0_t468[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t470 = FSM_fft_64_stage_6_0_t459;
    FSM_fft_64_stage_6_0_t470[FSM_fft_64_stage_6_0_t461 * 32 +: 32] = FSM_fft_64_stage_6_0_t469;
    FSM_fft_64_stage_6_0_t471 = 32'b00000000000000000000000000110111;
    FSM_fft_64_stage_6_0_t472 = FSM_fft_64_stage_6_0_t471[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t473 = 32'b00000000000000000000000000010111;
    FSM_fft_64_stage_6_0_t474 = FSM_fft_64_stage_6_0_t473[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t475 = i_data_in_real[FSM_fft_64_stage_6_0_t474 * 32 +: 32];
    FSM_fft_64_stage_6_0_t476 = 32'b00000000000000000000000000110111;
    FSM_fft_64_stage_6_0_t477 = FSM_fft_64_stage_6_0_t476[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t478 = i_data_in_real[FSM_fft_64_stage_6_0_t477 * 32 +: 32];
    FSM_fft_64_stage_6_0_t479 = FSM_fft_64_stage_6_0_t470;
    FSM_fft_64_stage_6_0_t479[FSM_fft_64_stage_6_0_t472 * 32 +: 32] = FSM_fft_64_stage_6_0_t475 - FSM_fft_64_stage_6_0_t478;
    FSM_fft_64_stage_6_0_t480 = 32'b00000000000000000000000000011000;
    FSM_fft_64_stage_6_0_t481 = FSM_fft_64_stage_6_0_t480[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t482 = 32'b00000000000000000000000000011000;
    FSM_fft_64_stage_6_0_t483 = FSM_fft_64_stage_6_0_t482[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t484 = i_data_in_real[FSM_fft_64_stage_6_0_t483 * 32 +: 32];
    FSM_fft_64_stage_6_0_t485 = 32'b00000000000000000000000000111000;
    FSM_fft_64_stage_6_0_t486 = FSM_fft_64_stage_6_0_t485[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t487 = i_data_in_real[FSM_fft_64_stage_6_0_t486 * 32 +: 32];
    FSM_fft_64_stage_6_0_t488 = FSM_fft_64_stage_6_0_t484 + FSM_fft_64_stage_6_0_t487;
    FSM_fft_64_stage_6_0_t489 = FSM_fft_64_stage_6_0_t488[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t490 = FSM_fft_64_stage_6_0_t479;
    FSM_fft_64_stage_6_0_t490[FSM_fft_64_stage_6_0_t481 * 32 +: 32] = FSM_fft_64_stage_6_0_t489;
    FSM_fft_64_stage_6_0_t491 = 32'b00000000000000000000000000111000;
    FSM_fft_64_stage_6_0_t492 = FSM_fft_64_stage_6_0_t491[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t493 = 32'b00000000000000000000000000011000;
    FSM_fft_64_stage_6_0_t494 = FSM_fft_64_stage_6_0_t493[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t495 = i_data_in_real[FSM_fft_64_stage_6_0_t494 * 32 +: 32];
    FSM_fft_64_stage_6_0_t496 = 32'b00000000000000000000000000111000;
    FSM_fft_64_stage_6_0_t497 = FSM_fft_64_stage_6_0_t496[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t498 = i_data_in_real[FSM_fft_64_stage_6_0_t497 * 32 +: 32];
    FSM_fft_64_stage_6_0_t499 = FSM_fft_64_stage_6_0_t490;
    FSM_fft_64_stage_6_0_t499[FSM_fft_64_stage_6_0_t492 * 32 +: 32] = FSM_fft_64_stage_6_0_t495 - FSM_fft_64_stage_6_0_t498;
    FSM_fft_64_stage_6_0_t500 = 32'b00000000000000000000000000011001;
    FSM_fft_64_stage_6_0_t501 = FSM_fft_64_stage_6_0_t500[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t502 = 32'b00000000000000000000000000011001;
    FSM_fft_64_stage_6_0_t503 = FSM_fft_64_stage_6_0_t502[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t504 = i_data_in_real[FSM_fft_64_stage_6_0_t503 * 32 +: 32];
    FSM_fft_64_stage_6_0_t505 = 32'b00000000000000000000000000111001;
    FSM_fft_64_stage_6_0_t506 = FSM_fft_64_stage_6_0_t505[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t507 = i_data_in_real[FSM_fft_64_stage_6_0_t506 * 32 +: 32];
    FSM_fft_64_stage_6_0_t508 = FSM_fft_64_stage_6_0_t504 + FSM_fft_64_stage_6_0_t507;
    FSM_fft_64_stage_6_0_t509 = FSM_fft_64_stage_6_0_t508[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t510 = FSM_fft_64_stage_6_0_t499;
    FSM_fft_64_stage_6_0_t510[FSM_fft_64_stage_6_0_t501 * 32 +: 32] = FSM_fft_64_stage_6_0_t509;
    FSM_fft_64_stage_6_0_t511 = 32'b00000000000000000000000000111001;
    FSM_fft_64_stage_6_0_t512 = FSM_fft_64_stage_6_0_t511[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t513 = 32'b00000000000000000000000000011001;
    FSM_fft_64_stage_6_0_t514 = FSM_fft_64_stage_6_0_t513[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t515 = i_data_in_real[FSM_fft_64_stage_6_0_t514 * 32 +: 32];
    FSM_fft_64_stage_6_0_t516 = 32'b00000000000000000000000000111001;
    FSM_fft_64_stage_6_0_t517 = FSM_fft_64_stage_6_0_t516[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t518 = i_data_in_real[FSM_fft_64_stage_6_0_t517 * 32 +: 32];
    FSM_fft_64_stage_6_0_t519 = FSM_fft_64_stage_6_0_t510;
    FSM_fft_64_stage_6_0_t519[FSM_fft_64_stage_6_0_t512 * 32 +: 32] = FSM_fft_64_stage_6_0_t515 - FSM_fft_64_stage_6_0_t518;
    FSM_fft_64_stage_6_0_t520 = 32'b00000000000000000000000000011010;
    FSM_fft_64_stage_6_0_t521 = FSM_fft_64_stage_6_0_t520[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t522 = 32'b00000000000000000000000000011010;
    FSM_fft_64_stage_6_0_t523 = FSM_fft_64_stage_6_0_t522[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t524 = i_data_in_real[FSM_fft_64_stage_6_0_t523 * 32 +: 32];
    FSM_fft_64_stage_6_0_t525 = 32'b00000000000000000000000000111010;
    FSM_fft_64_stage_6_0_t526 = FSM_fft_64_stage_6_0_t525[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t527 = i_data_in_real[FSM_fft_64_stage_6_0_t526 * 32 +: 32];
    FSM_fft_64_stage_6_0_t528 = FSM_fft_64_stage_6_0_t524 + FSM_fft_64_stage_6_0_t527;
    FSM_fft_64_stage_6_0_t529 = FSM_fft_64_stage_6_0_t528[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t530 = FSM_fft_64_stage_6_0_t519;
    FSM_fft_64_stage_6_0_t530[FSM_fft_64_stage_6_0_t521 * 32 +: 32] = FSM_fft_64_stage_6_0_t529;
    FSM_fft_64_stage_6_0_t531 = 32'b00000000000000000000000000111010;
    FSM_fft_64_stage_6_0_t532 = FSM_fft_64_stage_6_0_t531[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t533 = 32'b00000000000000000000000000011010;
    FSM_fft_64_stage_6_0_t534 = FSM_fft_64_stage_6_0_t533[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t535 = i_data_in_real[FSM_fft_64_stage_6_0_t534 * 32 +: 32];
    FSM_fft_64_stage_6_0_t536 = 32'b00000000000000000000000000111010;
    FSM_fft_64_stage_6_0_t537 = FSM_fft_64_stage_6_0_t536[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t538 = i_data_in_real[FSM_fft_64_stage_6_0_t537 * 32 +: 32];
    FSM_fft_64_stage_6_0_t539 = FSM_fft_64_stage_6_0_t530;
    FSM_fft_64_stage_6_0_t539[FSM_fft_64_stage_6_0_t532 * 32 +: 32] = FSM_fft_64_stage_6_0_t535 - FSM_fft_64_stage_6_0_t538;
    FSM_fft_64_stage_6_0_t540 = 32'b00000000000000000000000000011011;
    FSM_fft_64_stage_6_0_t541 = FSM_fft_64_stage_6_0_t540[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t542 = 32'b00000000000000000000000000011011;
    FSM_fft_64_stage_6_0_t543 = FSM_fft_64_stage_6_0_t542[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t544 = i_data_in_real[FSM_fft_64_stage_6_0_t543 * 32 +: 32];
    FSM_fft_64_stage_6_0_t545 = 32'b00000000000000000000000000111011;
    FSM_fft_64_stage_6_0_t546 = FSM_fft_64_stage_6_0_t545[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t547 = i_data_in_real[FSM_fft_64_stage_6_0_t546 * 32 +: 32];
    FSM_fft_64_stage_6_0_t548 = FSM_fft_64_stage_6_0_t544 + FSM_fft_64_stage_6_0_t547;
    FSM_fft_64_stage_6_0_t549 = FSM_fft_64_stage_6_0_t548[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t550 = FSM_fft_64_stage_6_0_t539;
    FSM_fft_64_stage_6_0_t550[FSM_fft_64_stage_6_0_t541 * 32 +: 32] = FSM_fft_64_stage_6_0_t549;
    FSM_fft_64_stage_6_0_t551 = 32'b00000000000000000000000000111011;
    FSM_fft_64_stage_6_0_t552 = FSM_fft_64_stage_6_0_t551[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t553 = 32'b00000000000000000000000000011011;
    FSM_fft_64_stage_6_0_t554 = FSM_fft_64_stage_6_0_t553[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t555 = i_data_in_real[FSM_fft_64_stage_6_0_t554 * 32 +: 32];
    FSM_fft_64_stage_6_0_t556 = 32'b00000000000000000000000000111011;
    FSM_fft_64_stage_6_0_t557 = FSM_fft_64_stage_6_0_t556[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t558 = i_data_in_real[FSM_fft_64_stage_6_0_t557 * 32 +: 32];
    FSM_fft_64_stage_6_0_t559 = FSM_fft_64_stage_6_0_t550;
    FSM_fft_64_stage_6_0_t559[FSM_fft_64_stage_6_0_t552 * 32 +: 32] = FSM_fft_64_stage_6_0_t555 - FSM_fft_64_stage_6_0_t558;
    FSM_fft_64_stage_6_0_t560 = 32'b00000000000000000000000000011100;
    FSM_fft_64_stage_6_0_t561 = FSM_fft_64_stage_6_0_t560[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t562 = 32'b00000000000000000000000000011100;
    FSM_fft_64_stage_6_0_t563 = FSM_fft_64_stage_6_0_t562[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t564 = i_data_in_real[FSM_fft_64_stage_6_0_t563 * 32 +: 32];
    FSM_fft_64_stage_6_0_t565 = 32'b00000000000000000000000000111100;
    FSM_fft_64_stage_6_0_t566 = FSM_fft_64_stage_6_0_t565[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t567 = i_data_in_real[FSM_fft_64_stage_6_0_t566 * 32 +: 32];
    FSM_fft_64_stage_6_0_t568 = FSM_fft_64_stage_6_0_t564 + FSM_fft_64_stage_6_0_t567;
    FSM_fft_64_stage_6_0_t569 = FSM_fft_64_stage_6_0_t568[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t570 = FSM_fft_64_stage_6_0_t559;
    FSM_fft_64_stage_6_0_t570[FSM_fft_64_stage_6_0_t561 * 32 +: 32] = FSM_fft_64_stage_6_0_t569;
    FSM_fft_64_stage_6_0_t571 = 32'b00000000000000000000000000111100;
    FSM_fft_64_stage_6_0_t572 = FSM_fft_64_stage_6_0_t571[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t573 = 32'b00000000000000000000000000011100;
    FSM_fft_64_stage_6_0_t574 = FSM_fft_64_stage_6_0_t573[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t575 = i_data_in_real[FSM_fft_64_stage_6_0_t574 * 32 +: 32];
    FSM_fft_64_stage_6_0_t576 = 32'b00000000000000000000000000111100;
    FSM_fft_64_stage_6_0_t577 = FSM_fft_64_stage_6_0_t576[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t578 = i_data_in_real[FSM_fft_64_stage_6_0_t577 * 32 +: 32];
    FSM_fft_64_stage_6_0_t579 = FSM_fft_64_stage_6_0_t570;
    FSM_fft_64_stage_6_0_t579[FSM_fft_64_stage_6_0_t572 * 32 +: 32] = FSM_fft_64_stage_6_0_t575 - FSM_fft_64_stage_6_0_t578;
    FSM_fft_64_stage_6_0_t580 = 32'b00000000000000000000000000011101;
    FSM_fft_64_stage_6_0_t581 = FSM_fft_64_stage_6_0_t580[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t582 = 32'b00000000000000000000000000011101;
    FSM_fft_64_stage_6_0_t583 = FSM_fft_64_stage_6_0_t582[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t584 = i_data_in_real[FSM_fft_64_stage_6_0_t583 * 32 +: 32];
    FSM_fft_64_stage_6_0_t585 = 32'b00000000000000000000000000111101;
    FSM_fft_64_stage_6_0_t586 = FSM_fft_64_stage_6_0_t585[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t587 = i_data_in_real[FSM_fft_64_stage_6_0_t586 * 32 +: 32];
    FSM_fft_64_stage_6_0_t588 = FSM_fft_64_stage_6_0_t584 + FSM_fft_64_stage_6_0_t587;
    FSM_fft_64_stage_6_0_t589 = FSM_fft_64_stage_6_0_t588[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t590 = FSM_fft_64_stage_6_0_t579;
    FSM_fft_64_stage_6_0_t590[FSM_fft_64_stage_6_0_t581 * 32 +: 32] = FSM_fft_64_stage_6_0_t589;
    FSM_fft_64_stage_6_0_t591 = 32'b00000000000000000000000000111101;
    FSM_fft_64_stage_6_0_t592 = FSM_fft_64_stage_6_0_t591[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t593 = 32'b00000000000000000000000000011101;
    FSM_fft_64_stage_6_0_t594 = FSM_fft_64_stage_6_0_t593[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t595 = i_data_in_real[FSM_fft_64_stage_6_0_t594 * 32 +: 32];
    FSM_fft_64_stage_6_0_t596 = 32'b00000000000000000000000000111101;
    FSM_fft_64_stage_6_0_t597 = FSM_fft_64_stage_6_0_t596[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t598 = i_data_in_real[FSM_fft_64_stage_6_0_t597 * 32 +: 32];
    FSM_fft_64_stage_6_0_t599 = FSM_fft_64_stage_6_0_t590;
    FSM_fft_64_stage_6_0_t599[FSM_fft_64_stage_6_0_t592 * 32 +: 32] = FSM_fft_64_stage_6_0_t595 - FSM_fft_64_stage_6_0_t598;
    FSM_fft_64_stage_6_0_t600 = 32'b00000000000000000000000000011110;
    FSM_fft_64_stage_6_0_t601 = FSM_fft_64_stage_6_0_t600[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t602 = 32'b00000000000000000000000000011110;
    FSM_fft_64_stage_6_0_t603 = FSM_fft_64_stage_6_0_t602[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t604 = i_data_in_real[FSM_fft_64_stage_6_0_t603 * 32 +: 32];
    FSM_fft_64_stage_6_0_t605 = 32'b00000000000000000000000000111110;
    FSM_fft_64_stage_6_0_t606 = FSM_fft_64_stage_6_0_t605[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t607 = i_data_in_real[FSM_fft_64_stage_6_0_t606 * 32 +: 32];
    FSM_fft_64_stage_6_0_t608 = FSM_fft_64_stage_6_0_t604 + FSM_fft_64_stage_6_0_t607;
    FSM_fft_64_stage_6_0_t609 = FSM_fft_64_stage_6_0_t608[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t610 = FSM_fft_64_stage_6_0_t599;
    FSM_fft_64_stage_6_0_t610[FSM_fft_64_stage_6_0_t601 * 32 +: 32] = FSM_fft_64_stage_6_0_t609;
    FSM_fft_64_stage_6_0_t611 = 32'b00000000000000000000000000111110;
    FSM_fft_64_stage_6_0_t612 = FSM_fft_64_stage_6_0_t611[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t613 = 32'b00000000000000000000000000011110;
    FSM_fft_64_stage_6_0_t614 = FSM_fft_64_stage_6_0_t613[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t615 = i_data_in_real[FSM_fft_64_stage_6_0_t614 * 32 +: 32];
    FSM_fft_64_stage_6_0_t616 = 32'b00000000000000000000000000111110;
    FSM_fft_64_stage_6_0_t617 = FSM_fft_64_stage_6_0_t616[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t618 = i_data_in_real[FSM_fft_64_stage_6_0_t617 * 32 +: 32];
    FSM_fft_64_stage_6_0_t619 = FSM_fft_64_stage_6_0_t610;
    FSM_fft_64_stage_6_0_t619[FSM_fft_64_stage_6_0_t612 * 32 +: 32] = FSM_fft_64_stage_6_0_t615 - FSM_fft_64_stage_6_0_t618;
    FSM_fft_64_stage_6_0_t620 = 32'b00000000000000000000000000011111;
    FSM_fft_64_stage_6_0_t621 = FSM_fft_64_stage_6_0_t620[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t622 = 32'b00000000000000000000000000011111;
    FSM_fft_64_stage_6_0_t623 = FSM_fft_64_stage_6_0_t622[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t624 = i_data_in_real[FSM_fft_64_stage_6_0_t623 * 32 +: 32];
    FSM_fft_64_stage_6_0_t625 = 32'b00000000000000000000000000111111;
    FSM_fft_64_stage_6_0_t626 = FSM_fft_64_stage_6_0_t625[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t627 = i_data_in_real[FSM_fft_64_stage_6_0_t626 * 32 +: 32];
    FSM_fft_64_stage_6_0_t628 = FSM_fft_64_stage_6_0_t624 + FSM_fft_64_stage_6_0_t627;
    FSM_fft_64_stage_6_0_t629 = FSM_fft_64_stage_6_0_t628[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t630 = FSM_fft_64_stage_6_0_t619;
    FSM_fft_64_stage_6_0_t630[FSM_fft_64_stage_6_0_t621 * 32 +: 32] = FSM_fft_64_stage_6_0_t629;
    FSM_fft_64_stage_6_0_t631 = 32'b00000000000000000000000000111111;
    FSM_fft_64_stage_6_0_t632 = FSM_fft_64_stage_6_0_t631[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t633 = 32'b00000000000000000000000000011111;
    FSM_fft_64_stage_6_0_t634 = FSM_fft_64_stage_6_0_t633[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t635 = i_data_in_real[FSM_fft_64_stage_6_0_t634 * 32 +: 32];
    FSM_fft_64_stage_6_0_t636 = 32'b00000000000000000000000000111111;
    FSM_fft_64_stage_6_0_t637 = FSM_fft_64_stage_6_0_t636[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t638 = i_data_in_real[FSM_fft_64_stage_6_0_t637 * 32 +: 32];
    FSM_fft_64_stage_6_0_t639 = FSM_fft_64_stage_6_0_t630;
    FSM_fft_64_stage_6_0_t639[FSM_fft_64_stage_6_0_t632 * 32 +: 32] = FSM_fft_64_stage_6_0_t635 - FSM_fft_64_stage_6_0_t638;
    FSM_fft_64_stage_6_0_t640 = 32'b0;
    FSM_fft_64_stage_6_0_t641 = FSM_fft_64_stage_6_0_t640[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t642 = 32'b0;
    FSM_fft_64_stage_6_0_t643 = FSM_fft_64_stage_6_0_t642[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t644 = i_data_in_imag[FSM_fft_64_stage_6_0_t643 * 32 +: 32];
    FSM_fft_64_stage_6_0_t645 = 32'b00000000000000000000000000100000;
    FSM_fft_64_stage_6_0_t646 = FSM_fft_64_stage_6_0_t645[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t647 = i_data_in_imag[FSM_fft_64_stage_6_0_t646 * 32 +: 32];
    FSM_fft_64_stage_6_0_t648 = FSM_fft_64_stage_6_0_t644 + FSM_fft_64_stage_6_0_t647;
    FSM_fft_64_stage_6_0_t649 = FSM_fft_64_stage_6_0_t648[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t650 = i_data_in_imag;
    FSM_fft_64_stage_6_0_t650[FSM_fft_64_stage_6_0_t641 * 32 +: 32] = FSM_fft_64_stage_6_0_t649;
    FSM_fft_64_stage_6_0_t651 = 32'b00000000000000000000000000100000;
    FSM_fft_64_stage_6_0_t652 = FSM_fft_64_stage_6_0_t651[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t653 = 32'b0;
    FSM_fft_64_stage_6_0_t654 = FSM_fft_64_stage_6_0_t653[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t655 = i_data_in_imag[FSM_fft_64_stage_6_0_t654 * 32 +: 32];
    FSM_fft_64_stage_6_0_t656 = 32'b00000000000000000000000000100000;
    FSM_fft_64_stage_6_0_t657 = FSM_fft_64_stage_6_0_t656[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t658 = i_data_in_imag[FSM_fft_64_stage_6_0_t657 * 32 +: 32];
    FSM_fft_64_stage_6_0_t659 = FSM_fft_64_stage_6_0_t650;
    FSM_fft_64_stage_6_0_t659[FSM_fft_64_stage_6_0_t652 * 32 +: 32] = FSM_fft_64_stage_6_0_t655 - FSM_fft_64_stage_6_0_t658;
    FSM_fft_64_stage_6_0_t660 = 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_6_0_t661 = FSM_fft_64_stage_6_0_t660[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t662 = 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_6_0_t663 = FSM_fft_64_stage_6_0_t662[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t664 = i_data_in_imag[FSM_fft_64_stage_6_0_t663 * 32 +: 32];
    FSM_fft_64_stage_6_0_t665 = 32'b00000000000000000000000000100001;
    FSM_fft_64_stage_6_0_t666 = FSM_fft_64_stage_6_0_t665[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t667 = i_data_in_imag[FSM_fft_64_stage_6_0_t666 * 32 +: 32];
    FSM_fft_64_stage_6_0_t668 = FSM_fft_64_stage_6_0_t664 + FSM_fft_64_stage_6_0_t667;
    FSM_fft_64_stage_6_0_t669 = FSM_fft_64_stage_6_0_t668[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t670 = FSM_fft_64_stage_6_0_t659;
    FSM_fft_64_stage_6_0_t670[FSM_fft_64_stage_6_0_t661 * 32 +: 32] = FSM_fft_64_stage_6_0_t669;
    FSM_fft_64_stage_6_0_t671 = 32'b00000000000000000000000000100001;
    FSM_fft_64_stage_6_0_t672 = FSM_fft_64_stage_6_0_t671[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t673 = 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_6_0_t674 = FSM_fft_64_stage_6_0_t673[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t675 = i_data_in_imag[FSM_fft_64_stage_6_0_t674 * 32 +: 32];
    FSM_fft_64_stage_6_0_t676 = 32'b00000000000000000000000000100001;
    FSM_fft_64_stage_6_0_t677 = FSM_fft_64_stage_6_0_t676[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t678 = i_data_in_imag[FSM_fft_64_stage_6_0_t677 * 32 +: 32];
    FSM_fft_64_stage_6_0_t679 = FSM_fft_64_stage_6_0_t670;
    FSM_fft_64_stage_6_0_t679[FSM_fft_64_stage_6_0_t672 * 32 +: 32] = FSM_fft_64_stage_6_0_t675 - FSM_fft_64_stage_6_0_t678;
    FSM_fft_64_stage_6_0_t680 = 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_6_0_t681 = FSM_fft_64_stage_6_0_t680[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t682 = 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_6_0_t683 = FSM_fft_64_stage_6_0_t682[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t684 = i_data_in_imag[FSM_fft_64_stage_6_0_t683 * 32 +: 32];
    FSM_fft_64_stage_6_0_t685 = 32'b00000000000000000000000000100010;
    FSM_fft_64_stage_6_0_t686 = FSM_fft_64_stage_6_0_t685[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t687 = i_data_in_imag[FSM_fft_64_stage_6_0_t686 * 32 +: 32];
    FSM_fft_64_stage_6_0_t688 = FSM_fft_64_stage_6_0_t684 + FSM_fft_64_stage_6_0_t687;
    FSM_fft_64_stage_6_0_t689 = FSM_fft_64_stage_6_0_t688[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t690 = FSM_fft_64_stage_6_0_t679;
    FSM_fft_64_stage_6_0_t690[FSM_fft_64_stage_6_0_t681 * 32 +: 32] = FSM_fft_64_stage_6_0_t689;
    FSM_fft_64_stage_6_0_t691 = 32'b00000000000000000000000000100010;
    FSM_fft_64_stage_6_0_t692 = FSM_fft_64_stage_6_0_t691[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t693 = 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_6_0_t694 = FSM_fft_64_stage_6_0_t693[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t695 = i_data_in_imag[FSM_fft_64_stage_6_0_t694 * 32 +: 32];
    FSM_fft_64_stage_6_0_t696 = 32'b00000000000000000000000000100010;
    FSM_fft_64_stage_6_0_t697 = FSM_fft_64_stage_6_0_t696[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t698 = i_data_in_imag[FSM_fft_64_stage_6_0_t697 * 32 +: 32];
    FSM_fft_64_stage_6_0_t699 = FSM_fft_64_stage_6_0_t690;
    FSM_fft_64_stage_6_0_t699[FSM_fft_64_stage_6_0_t692 * 32 +: 32] = FSM_fft_64_stage_6_0_t695 - FSM_fft_64_stage_6_0_t698;
    FSM_fft_64_stage_6_0_t700 = 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_6_0_t701 = FSM_fft_64_stage_6_0_t700[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t702 = 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_6_0_t703 = FSM_fft_64_stage_6_0_t702[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t704 = i_data_in_imag[FSM_fft_64_stage_6_0_t703 * 32 +: 32];
    FSM_fft_64_stage_6_0_t705 = 32'b00000000000000000000000000100011;
    FSM_fft_64_stage_6_0_t706 = FSM_fft_64_stage_6_0_t705[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t707 = i_data_in_imag[FSM_fft_64_stage_6_0_t706 * 32 +: 32];
    FSM_fft_64_stage_6_0_t708 = FSM_fft_64_stage_6_0_t704 + FSM_fft_64_stage_6_0_t707;
    FSM_fft_64_stage_6_0_t709 = FSM_fft_64_stage_6_0_t708[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t710 = FSM_fft_64_stage_6_0_t699;
    FSM_fft_64_stage_6_0_t710[FSM_fft_64_stage_6_0_t701 * 32 +: 32] = FSM_fft_64_stage_6_0_t709;
    FSM_fft_64_stage_6_0_t711 = 32'b00000000000000000000000000100011;
    FSM_fft_64_stage_6_0_t712 = FSM_fft_64_stage_6_0_t711[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t713 = 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_6_0_t714 = FSM_fft_64_stage_6_0_t713[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t715 = i_data_in_imag[FSM_fft_64_stage_6_0_t714 * 32 +: 32];
    FSM_fft_64_stage_6_0_t716 = 32'b00000000000000000000000000100011;
    FSM_fft_64_stage_6_0_t717 = FSM_fft_64_stage_6_0_t716[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t718 = i_data_in_imag[FSM_fft_64_stage_6_0_t717 * 32 +: 32];
    FSM_fft_64_stage_6_0_t719 = FSM_fft_64_stage_6_0_t710;
    FSM_fft_64_stage_6_0_t719[FSM_fft_64_stage_6_0_t712 * 32 +: 32] = FSM_fft_64_stage_6_0_t715 - FSM_fft_64_stage_6_0_t718;
    FSM_fft_64_stage_6_0_t720 = 32'b00000000000000000000000000000100;
    FSM_fft_64_stage_6_0_t721 = FSM_fft_64_stage_6_0_t720[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t722 = 32'b00000000000000000000000000000100;
    FSM_fft_64_stage_6_0_t723 = FSM_fft_64_stage_6_0_t722[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t724 = i_data_in_imag[FSM_fft_64_stage_6_0_t723 * 32 +: 32];
    FSM_fft_64_stage_6_0_t725 = 32'b00000000000000000000000000100100;
    FSM_fft_64_stage_6_0_t726 = FSM_fft_64_stage_6_0_t725[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t727 = i_data_in_imag[FSM_fft_64_stage_6_0_t726 * 32 +: 32];
    FSM_fft_64_stage_6_0_t728 = FSM_fft_64_stage_6_0_t724 + FSM_fft_64_stage_6_0_t727;
    FSM_fft_64_stage_6_0_t729 = FSM_fft_64_stage_6_0_t728[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t730 = FSM_fft_64_stage_6_0_t719;
    FSM_fft_64_stage_6_0_t730[FSM_fft_64_stage_6_0_t721 * 32 +: 32] = FSM_fft_64_stage_6_0_t729;
    FSM_fft_64_stage_6_0_t731 = 32'b00000000000000000000000000100100;
    FSM_fft_64_stage_6_0_t732 = FSM_fft_64_stage_6_0_t731[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t733 = 32'b00000000000000000000000000000100;
    FSM_fft_64_stage_6_0_t734 = FSM_fft_64_stage_6_0_t733[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t735 = i_data_in_imag[FSM_fft_64_stage_6_0_t734 * 32 +: 32];
    FSM_fft_64_stage_6_0_t736 = 32'b00000000000000000000000000100100;
    FSM_fft_64_stage_6_0_t737 = FSM_fft_64_stage_6_0_t736[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t738 = i_data_in_imag[FSM_fft_64_stage_6_0_t737 * 32 +: 32];
    FSM_fft_64_stage_6_0_t739 = FSM_fft_64_stage_6_0_t730;
    FSM_fft_64_stage_6_0_t739[FSM_fft_64_stage_6_0_t732 * 32 +: 32] = FSM_fft_64_stage_6_0_t735 - FSM_fft_64_stage_6_0_t738;
    FSM_fft_64_stage_6_0_t740 = 32'b00000000000000000000000000000101;
    FSM_fft_64_stage_6_0_t741 = FSM_fft_64_stage_6_0_t740[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t742 = 32'b00000000000000000000000000000101;
    FSM_fft_64_stage_6_0_t743 = FSM_fft_64_stage_6_0_t742[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t744 = i_data_in_imag[FSM_fft_64_stage_6_0_t743 * 32 +: 32];
    FSM_fft_64_stage_6_0_t745 = 32'b00000000000000000000000000100101;
    FSM_fft_64_stage_6_0_t746 = FSM_fft_64_stage_6_0_t745[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t747 = i_data_in_imag[FSM_fft_64_stage_6_0_t746 * 32 +: 32];
    FSM_fft_64_stage_6_0_t748 = FSM_fft_64_stage_6_0_t744 + FSM_fft_64_stage_6_0_t747;
    FSM_fft_64_stage_6_0_t749 = FSM_fft_64_stage_6_0_t748[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t750 = FSM_fft_64_stage_6_0_t739;
    FSM_fft_64_stage_6_0_t750[FSM_fft_64_stage_6_0_t741 * 32 +: 32] = FSM_fft_64_stage_6_0_t749;
    FSM_fft_64_stage_6_0_t751 = 32'b00000000000000000000000000100101;
    FSM_fft_64_stage_6_0_t752 = FSM_fft_64_stage_6_0_t751[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t753 = 32'b00000000000000000000000000000101;
    FSM_fft_64_stage_6_0_t754 = FSM_fft_64_stage_6_0_t753[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t755 = i_data_in_imag[FSM_fft_64_stage_6_0_t754 * 32 +: 32];
    FSM_fft_64_stage_6_0_t756 = 32'b00000000000000000000000000100101;
    FSM_fft_64_stage_6_0_t757 = FSM_fft_64_stage_6_0_t756[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t758 = i_data_in_imag[FSM_fft_64_stage_6_0_t757 * 32 +: 32];
    FSM_fft_64_stage_6_0_t759 = FSM_fft_64_stage_6_0_t750;
    FSM_fft_64_stage_6_0_t759[FSM_fft_64_stage_6_0_t752 * 32 +: 32] = FSM_fft_64_stage_6_0_t755 - FSM_fft_64_stage_6_0_t758;
    FSM_fft_64_stage_6_0_t760 = 32'b00000000000000000000000000000110;
    FSM_fft_64_stage_6_0_t761 = FSM_fft_64_stage_6_0_t760[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t762 = 32'b00000000000000000000000000000110;
    FSM_fft_64_stage_6_0_t763 = FSM_fft_64_stage_6_0_t762[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t764 = i_data_in_imag[FSM_fft_64_stage_6_0_t763 * 32 +: 32];
    FSM_fft_64_stage_6_0_t765 = 32'b00000000000000000000000000100110;
    FSM_fft_64_stage_6_0_t766 = FSM_fft_64_stage_6_0_t765[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t767 = i_data_in_imag[FSM_fft_64_stage_6_0_t766 * 32 +: 32];
    FSM_fft_64_stage_6_0_t768 = FSM_fft_64_stage_6_0_t764 + FSM_fft_64_stage_6_0_t767;
    FSM_fft_64_stage_6_0_t769 = FSM_fft_64_stage_6_0_t768[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t770 = FSM_fft_64_stage_6_0_t759;
    FSM_fft_64_stage_6_0_t770[FSM_fft_64_stage_6_0_t761 * 32 +: 32] = FSM_fft_64_stage_6_0_t769;
    FSM_fft_64_stage_6_0_t771 = 32'b00000000000000000000000000100110;
    FSM_fft_64_stage_6_0_t772 = FSM_fft_64_stage_6_0_t771[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t773 = 32'b00000000000000000000000000000110;
    FSM_fft_64_stage_6_0_t774 = FSM_fft_64_stage_6_0_t773[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t775 = i_data_in_imag[FSM_fft_64_stage_6_0_t774 * 32 +: 32];
    FSM_fft_64_stage_6_0_t776 = 32'b00000000000000000000000000100110;
    FSM_fft_64_stage_6_0_t777 = FSM_fft_64_stage_6_0_t776[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t778 = i_data_in_imag[FSM_fft_64_stage_6_0_t777 * 32 +: 32];
    FSM_fft_64_stage_6_0_t779 = FSM_fft_64_stage_6_0_t770;
    FSM_fft_64_stage_6_0_t779[FSM_fft_64_stage_6_0_t772 * 32 +: 32] = FSM_fft_64_stage_6_0_t775 - FSM_fft_64_stage_6_0_t778;
    FSM_fft_64_stage_6_0_t780 = 32'b00000000000000000000000000000111;
    FSM_fft_64_stage_6_0_t781 = FSM_fft_64_stage_6_0_t780[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t782 = 32'b00000000000000000000000000000111;
    FSM_fft_64_stage_6_0_t783 = FSM_fft_64_stage_6_0_t782[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t784 = i_data_in_imag[FSM_fft_64_stage_6_0_t783 * 32 +: 32];
    FSM_fft_64_stage_6_0_t785 = 32'b00000000000000000000000000100111;
    FSM_fft_64_stage_6_0_t786 = FSM_fft_64_stage_6_0_t785[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t787 = i_data_in_imag[FSM_fft_64_stage_6_0_t786 * 32 +: 32];
    FSM_fft_64_stage_6_0_t788 = FSM_fft_64_stage_6_0_t784 + FSM_fft_64_stage_6_0_t787;
    FSM_fft_64_stage_6_0_t789 = FSM_fft_64_stage_6_0_t788[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t790 = FSM_fft_64_stage_6_0_t779;
    FSM_fft_64_stage_6_0_t790[FSM_fft_64_stage_6_0_t781 * 32 +: 32] = FSM_fft_64_stage_6_0_t789;
    FSM_fft_64_stage_6_0_t791 = 32'b00000000000000000000000000100111;
    FSM_fft_64_stage_6_0_t792 = FSM_fft_64_stage_6_0_t791[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t793 = 32'b00000000000000000000000000000111;
    FSM_fft_64_stage_6_0_t794 = FSM_fft_64_stage_6_0_t793[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t795 = i_data_in_imag[FSM_fft_64_stage_6_0_t794 * 32 +: 32];
    FSM_fft_64_stage_6_0_t796 = 32'b00000000000000000000000000100111;
    FSM_fft_64_stage_6_0_t797 = FSM_fft_64_stage_6_0_t796[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t798 = i_data_in_imag[FSM_fft_64_stage_6_0_t797 * 32 +: 32];
    FSM_fft_64_stage_6_0_t799 = FSM_fft_64_stage_6_0_t790;
    FSM_fft_64_stage_6_0_t799[FSM_fft_64_stage_6_0_t792 * 32 +: 32] = FSM_fft_64_stage_6_0_t795 - FSM_fft_64_stage_6_0_t798;
    FSM_fft_64_stage_6_0_t800 = 32'b00000000000000000000000000001000;
    FSM_fft_64_stage_6_0_t801 = FSM_fft_64_stage_6_0_t800[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t802 = 32'b00000000000000000000000000001000;
    FSM_fft_64_stage_6_0_t803 = FSM_fft_64_stage_6_0_t802[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t804 = i_data_in_imag[FSM_fft_64_stage_6_0_t803 * 32 +: 32];
    FSM_fft_64_stage_6_0_t805 = 32'b00000000000000000000000000101000;
    FSM_fft_64_stage_6_0_t806 = FSM_fft_64_stage_6_0_t805[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t807 = i_data_in_imag[FSM_fft_64_stage_6_0_t806 * 32 +: 32];
    FSM_fft_64_stage_6_0_t808 = FSM_fft_64_stage_6_0_t804 + FSM_fft_64_stage_6_0_t807;
    FSM_fft_64_stage_6_0_t809 = FSM_fft_64_stage_6_0_t808[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t810 = FSM_fft_64_stage_6_0_t799;
    FSM_fft_64_stage_6_0_t810[FSM_fft_64_stage_6_0_t801 * 32 +: 32] = FSM_fft_64_stage_6_0_t809;
    FSM_fft_64_stage_6_0_t811 = 32'b00000000000000000000000000101000;
    FSM_fft_64_stage_6_0_t812 = FSM_fft_64_stage_6_0_t811[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t813 = 32'b00000000000000000000000000001000;
    FSM_fft_64_stage_6_0_t814 = FSM_fft_64_stage_6_0_t813[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t815 = i_data_in_imag[FSM_fft_64_stage_6_0_t814 * 32 +: 32];
    FSM_fft_64_stage_6_0_t816 = 32'b00000000000000000000000000101000;
    FSM_fft_64_stage_6_0_t817 = FSM_fft_64_stage_6_0_t816[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t818 = i_data_in_imag[FSM_fft_64_stage_6_0_t817 * 32 +: 32];
    FSM_fft_64_stage_6_0_t819 = FSM_fft_64_stage_6_0_t810;
    FSM_fft_64_stage_6_0_t819[FSM_fft_64_stage_6_0_t812 * 32 +: 32] = FSM_fft_64_stage_6_0_t815 - FSM_fft_64_stage_6_0_t818;
    FSM_fft_64_stage_6_0_t820 = 32'b00000000000000000000000000001001;
    FSM_fft_64_stage_6_0_t821 = FSM_fft_64_stage_6_0_t820[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t822 = 32'b00000000000000000000000000001001;
    FSM_fft_64_stage_6_0_t823 = FSM_fft_64_stage_6_0_t822[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t824 = i_data_in_imag[FSM_fft_64_stage_6_0_t823 * 32 +: 32];
    FSM_fft_64_stage_6_0_t825 = 32'b00000000000000000000000000101001;
    FSM_fft_64_stage_6_0_t826 = FSM_fft_64_stage_6_0_t825[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t827 = i_data_in_imag[FSM_fft_64_stage_6_0_t826 * 32 +: 32];
    FSM_fft_64_stage_6_0_t828 = FSM_fft_64_stage_6_0_t824 + FSM_fft_64_stage_6_0_t827;
    FSM_fft_64_stage_6_0_t829 = FSM_fft_64_stage_6_0_t828[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t830 = FSM_fft_64_stage_6_0_t819;
    FSM_fft_64_stage_6_0_t830[FSM_fft_64_stage_6_0_t821 * 32 +: 32] = FSM_fft_64_stage_6_0_t829;
    FSM_fft_64_stage_6_0_t831 = 32'b00000000000000000000000000101001;
    FSM_fft_64_stage_6_0_t832 = FSM_fft_64_stage_6_0_t831[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t833 = 32'b00000000000000000000000000001001;
    FSM_fft_64_stage_6_0_t834 = FSM_fft_64_stage_6_0_t833[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t835 = i_data_in_imag[FSM_fft_64_stage_6_0_t834 * 32 +: 32];
    FSM_fft_64_stage_6_0_t836 = 32'b00000000000000000000000000101001;
    FSM_fft_64_stage_6_0_t837 = FSM_fft_64_stage_6_0_t836[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t838 = i_data_in_imag[FSM_fft_64_stage_6_0_t837 * 32 +: 32];
    FSM_fft_64_stage_6_0_t839 = FSM_fft_64_stage_6_0_t830;
    FSM_fft_64_stage_6_0_t839[FSM_fft_64_stage_6_0_t832 * 32 +: 32] = FSM_fft_64_stage_6_0_t835 - FSM_fft_64_stage_6_0_t838;
    FSM_fft_64_stage_6_0_t840 = 32'b00000000000000000000000000001010;
    FSM_fft_64_stage_6_0_t841 = FSM_fft_64_stage_6_0_t840[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t842 = 32'b00000000000000000000000000001010;
    FSM_fft_64_stage_6_0_t843 = FSM_fft_64_stage_6_0_t842[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t844 = i_data_in_imag[FSM_fft_64_stage_6_0_t843 * 32 +: 32];
    FSM_fft_64_stage_6_0_t845 = 32'b00000000000000000000000000101010;
    FSM_fft_64_stage_6_0_t846 = FSM_fft_64_stage_6_0_t845[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t847 = i_data_in_imag[FSM_fft_64_stage_6_0_t846 * 32 +: 32];
    FSM_fft_64_stage_6_0_t848 = FSM_fft_64_stage_6_0_t844 + FSM_fft_64_stage_6_0_t847;
    FSM_fft_64_stage_6_0_t849 = FSM_fft_64_stage_6_0_t848[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t850 = FSM_fft_64_stage_6_0_t839;
    FSM_fft_64_stage_6_0_t850[FSM_fft_64_stage_6_0_t841 * 32 +: 32] = FSM_fft_64_stage_6_0_t849;
    FSM_fft_64_stage_6_0_t851 = 32'b00000000000000000000000000101010;
    FSM_fft_64_stage_6_0_t852 = FSM_fft_64_stage_6_0_t851[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t853 = 32'b00000000000000000000000000001010;
    FSM_fft_64_stage_6_0_t854 = FSM_fft_64_stage_6_0_t853[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t855 = i_data_in_imag[FSM_fft_64_stage_6_0_t854 * 32 +: 32];
    FSM_fft_64_stage_6_0_t856 = 32'b00000000000000000000000000101010;
    FSM_fft_64_stage_6_0_t857 = FSM_fft_64_stage_6_0_t856[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t858 = i_data_in_imag[FSM_fft_64_stage_6_0_t857 * 32 +: 32];
    FSM_fft_64_stage_6_0_t859 = FSM_fft_64_stage_6_0_t850;
    FSM_fft_64_stage_6_0_t859[FSM_fft_64_stage_6_0_t852 * 32 +: 32] = FSM_fft_64_stage_6_0_t855 - FSM_fft_64_stage_6_0_t858;
    FSM_fft_64_stage_6_0_t860 = 32'b00000000000000000000000000001011;
    FSM_fft_64_stage_6_0_t861 = FSM_fft_64_stage_6_0_t860[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t862 = 32'b00000000000000000000000000001011;
    FSM_fft_64_stage_6_0_t863 = FSM_fft_64_stage_6_0_t862[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t864 = i_data_in_imag[FSM_fft_64_stage_6_0_t863 * 32 +: 32];
    FSM_fft_64_stage_6_0_t865 = 32'b00000000000000000000000000101011;
    FSM_fft_64_stage_6_0_t866 = FSM_fft_64_stage_6_0_t865[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t867 = i_data_in_imag[FSM_fft_64_stage_6_0_t866 * 32 +: 32];
    FSM_fft_64_stage_6_0_t868 = FSM_fft_64_stage_6_0_t864 + FSM_fft_64_stage_6_0_t867;
    FSM_fft_64_stage_6_0_t869 = FSM_fft_64_stage_6_0_t868[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t870 = FSM_fft_64_stage_6_0_t859;
    FSM_fft_64_stage_6_0_t870[FSM_fft_64_stage_6_0_t861 * 32 +: 32] = FSM_fft_64_stage_6_0_t869;
    FSM_fft_64_stage_6_0_t871 = 32'b00000000000000000000000000101011;
    FSM_fft_64_stage_6_0_t872 = FSM_fft_64_stage_6_0_t871[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t873 = 32'b00000000000000000000000000001011;
    FSM_fft_64_stage_6_0_t874 = FSM_fft_64_stage_6_0_t873[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t875 = i_data_in_imag[FSM_fft_64_stage_6_0_t874 * 32 +: 32];
    FSM_fft_64_stage_6_0_t876 = 32'b00000000000000000000000000101011;
    FSM_fft_64_stage_6_0_t877 = FSM_fft_64_stage_6_0_t876[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t878 = i_data_in_imag[FSM_fft_64_stage_6_0_t877 * 32 +: 32];
    FSM_fft_64_stage_6_0_t879 = FSM_fft_64_stage_6_0_t870;
    FSM_fft_64_stage_6_0_t879[FSM_fft_64_stage_6_0_t872 * 32 +: 32] = FSM_fft_64_stage_6_0_t875 - FSM_fft_64_stage_6_0_t878;
    FSM_fft_64_stage_6_0_t880 = 32'b00000000000000000000000000001100;
    FSM_fft_64_stage_6_0_t881 = FSM_fft_64_stage_6_0_t880[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t882 = 32'b00000000000000000000000000001100;
    FSM_fft_64_stage_6_0_t883 = FSM_fft_64_stage_6_0_t882[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t884 = i_data_in_imag[FSM_fft_64_stage_6_0_t883 * 32 +: 32];
    FSM_fft_64_stage_6_0_t885 = 32'b00000000000000000000000000101100;
    FSM_fft_64_stage_6_0_t886 = FSM_fft_64_stage_6_0_t885[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t887 = i_data_in_imag[FSM_fft_64_stage_6_0_t886 * 32 +: 32];
    FSM_fft_64_stage_6_0_t888 = FSM_fft_64_stage_6_0_t884 + FSM_fft_64_stage_6_0_t887;
    FSM_fft_64_stage_6_0_t889 = FSM_fft_64_stage_6_0_t888[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t890 = FSM_fft_64_stage_6_0_t879;
    FSM_fft_64_stage_6_0_t890[FSM_fft_64_stage_6_0_t881 * 32 +: 32] = FSM_fft_64_stage_6_0_t889;
    FSM_fft_64_stage_6_0_t891 = 32'b00000000000000000000000000101100;
    FSM_fft_64_stage_6_0_t892 = FSM_fft_64_stage_6_0_t891[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t893 = 32'b00000000000000000000000000001100;
    FSM_fft_64_stage_6_0_t894 = FSM_fft_64_stage_6_0_t893[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t895 = i_data_in_imag[FSM_fft_64_stage_6_0_t894 * 32 +: 32];
    FSM_fft_64_stage_6_0_t896 = 32'b00000000000000000000000000101100;
    FSM_fft_64_stage_6_0_t897 = FSM_fft_64_stage_6_0_t896[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t898 = i_data_in_imag[FSM_fft_64_stage_6_0_t897 * 32 +: 32];
    FSM_fft_64_stage_6_0_t899 = FSM_fft_64_stage_6_0_t890;
    FSM_fft_64_stage_6_0_t899[FSM_fft_64_stage_6_0_t892 * 32 +: 32] = FSM_fft_64_stage_6_0_t895 - FSM_fft_64_stage_6_0_t898;
    FSM_fft_64_stage_6_0_t900 = 32'b00000000000000000000000000001101;
    FSM_fft_64_stage_6_0_t901 = FSM_fft_64_stage_6_0_t900[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t902 = 32'b00000000000000000000000000001101;
    FSM_fft_64_stage_6_0_t903 = FSM_fft_64_stage_6_0_t902[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t904 = i_data_in_imag[FSM_fft_64_stage_6_0_t903 * 32 +: 32];
    FSM_fft_64_stage_6_0_t905 = 32'b00000000000000000000000000101101;
    FSM_fft_64_stage_6_0_t906 = FSM_fft_64_stage_6_0_t905[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t907 = i_data_in_imag[FSM_fft_64_stage_6_0_t906 * 32 +: 32];
    FSM_fft_64_stage_6_0_t908 = FSM_fft_64_stage_6_0_t904 + FSM_fft_64_stage_6_0_t907;
    FSM_fft_64_stage_6_0_t909 = FSM_fft_64_stage_6_0_t908[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t910 = FSM_fft_64_stage_6_0_t899;
    FSM_fft_64_stage_6_0_t910[FSM_fft_64_stage_6_0_t901 * 32 +: 32] = FSM_fft_64_stage_6_0_t909;
    FSM_fft_64_stage_6_0_t911 = 32'b00000000000000000000000000101101;
    FSM_fft_64_stage_6_0_t912 = FSM_fft_64_stage_6_0_t911[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t913 = 32'b00000000000000000000000000001101;
    FSM_fft_64_stage_6_0_t914 = FSM_fft_64_stage_6_0_t913[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t915 = i_data_in_imag[FSM_fft_64_stage_6_0_t914 * 32 +: 32];
    FSM_fft_64_stage_6_0_t916 = 32'b00000000000000000000000000101101;
    FSM_fft_64_stage_6_0_t917 = FSM_fft_64_stage_6_0_t916[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t918 = i_data_in_imag[FSM_fft_64_stage_6_0_t917 * 32 +: 32];
    FSM_fft_64_stage_6_0_t919 = FSM_fft_64_stage_6_0_t910;
    FSM_fft_64_stage_6_0_t919[FSM_fft_64_stage_6_0_t912 * 32 +: 32] = FSM_fft_64_stage_6_0_t915 - FSM_fft_64_stage_6_0_t918;
    FSM_fft_64_stage_6_0_t920 = 32'b00000000000000000000000000001110;
    FSM_fft_64_stage_6_0_t921 = FSM_fft_64_stage_6_0_t920[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t922 = 32'b00000000000000000000000000001110;
    FSM_fft_64_stage_6_0_t923 = FSM_fft_64_stage_6_0_t922[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t924 = i_data_in_imag[FSM_fft_64_stage_6_0_t923 * 32 +: 32];
    FSM_fft_64_stage_6_0_t925 = 32'b00000000000000000000000000101110;
    FSM_fft_64_stage_6_0_t926 = FSM_fft_64_stage_6_0_t925[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t927 = i_data_in_imag[FSM_fft_64_stage_6_0_t926 * 32 +: 32];
    FSM_fft_64_stage_6_0_t928 = FSM_fft_64_stage_6_0_t924 + FSM_fft_64_stage_6_0_t927;
    FSM_fft_64_stage_6_0_t929 = FSM_fft_64_stage_6_0_t928[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t930 = FSM_fft_64_stage_6_0_t919;
    FSM_fft_64_stage_6_0_t930[FSM_fft_64_stage_6_0_t921 * 32 +: 32] = FSM_fft_64_stage_6_0_t929;
    FSM_fft_64_stage_6_0_t931 = 32'b00000000000000000000000000101110;
    FSM_fft_64_stage_6_0_t932 = FSM_fft_64_stage_6_0_t931[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t933 = 32'b00000000000000000000000000001110;
    FSM_fft_64_stage_6_0_t934 = FSM_fft_64_stage_6_0_t933[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t935 = i_data_in_imag[FSM_fft_64_stage_6_0_t934 * 32 +: 32];
    FSM_fft_64_stage_6_0_t936 = 32'b00000000000000000000000000101110;
    FSM_fft_64_stage_6_0_t937 = FSM_fft_64_stage_6_0_t936[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t938 = i_data_in_imag[FSM_fft_64_stage_6_0_t937 * 32 +: 32];
    FSM_fft_64_stage_6_0_t939 = FSM_fft_64_stage_6_0_t930;
    FSM_fft_64_stage_6_0_t939[FSM_fft_64_stage_6_0_t932 * 32 +: 32] = FSM_fft_64_stage_6_0_t935 - FSM_fft_64_stage_6_0_t938;
    FSM_fft_64_stage_6_0_t940 = 32'b00000000000000000000000000001111;
    FSM_fft_64_stage_6_0_t941 = FSM_fft_64_stage_6_0_t940[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t942 = 32'b00000000000000000000000000001111;
    FSM_fft_64_stage_6_0_t943 = FSM_fft_64_stage_6_0_t942[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t944 = i_data_in_imag[FSM_fft_64_stage_6_0_t943 * 32 +: 32];
    FSM_fft_64_stage_6_0_t945 = 32'b00000000000000000000000000101111;
    FSM_fft_64_stage_6_0_t946 = FSM_fft_64_stage_6_0_t945[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t947 = i_data_in_imag[FSM_fft_64_stage_6_0_t946 * 32 +: 32];
    FSM_fft_64_stage_6_0_t948 = FSM_fft_64_stage_6_0_t944 + FSM_fft_64_stage_6_0_t947;
    FSM_fft_64_stage_6_0_t949 = FSM_fft_64_stage_6_0_t948[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t950 = FSM_fft_64_stage_6_0_t939;
    FSM_fft_64_stage_6_0_t950[FSM_fft_64_stage_6_0_t941 * 32 +: 32] = FSM_fft_64_stage_6_0_t949;
    FSM_fft_64_stage_6_0_t951 = 32'b00000000000000000000000000101111;
    FSM_fft_64_stage_6_0_t952 = FSM_fft_64_stage_6_0_t951[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t953 = 32'b00000000000000000000000000001111;
    FSM_fft_64_stage_6_0_t954 = FSM_fft_64_stage_6_0_t953[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t955 = i_data_in_imag[FSM_fft_64_stage_6_0_t954 * 32 +: 32];
    FSM_fft_64_stage_6_0_t956 = 32'b00000000000000000000000000101111;
    FSM_fft_64_stage_6_0_t957 = FSM_fft_64_stage_6_0_t956[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t958 = i_data_in_imag[FSM_fft_64_stage_6_0_t957 * 32 +: 32];
    FSM_fft_64_stage_6_0_t959 = FSM_fft_64_stage_6_0_t950;
    FSM_fft_64_stage_6_0_t959[FSM_fft_64_stage_6_0_t952 * 32 +: 32] = FSM_fft_64_stage_6_0_t955 - FSM_fft_64_stage_6_0_t958;
    FSM_fft_64_stage_6_0_t960 = 32'b00000000000000000000000000010000;
    FSM_fft_64_stage_6_0_t961 = FSM_fft_64_stage_6_0_t960[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t962 = 32'b00000000000000000000000000010000;
    FSM_fft_64_stage_6_0_t963 = FSM_fft_64_stage_6_0_t962[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t964 = i_data_in_imag[FSM_fft_64_stage_6_0_t963 * 32 +: 32];
    FSM_fft_64_stage_6_0_t965 = 32'b00000000000000000000000000110000;
    FSM_fft_64_stage_6_0_t966 = FSM_fft_64_stage_6_0_t965[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t967 = i_data_in_imag[FSM_fft_64_stage_6_0_t966 * 32 +: 32];
    FSM_fft_64_stage_6_0_t968 = FSM_fft_64_stage_6_0_t964 + FSM_fft_64_stage_6_0_t967;
    FSM_fft_64_stage_6_0_t969 = FSM_fft_64_stage_6_0_t968[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t970 = FSM_fft_64_stage_6_0_t959;
    FSM_fft_64_stage_6_0_t970[FSM_fft_64_stage_6_0_t961 * 32 +: 32] = FSM_fft_64_stage_6_0_t969;
    FSM_fft_64_stage_6_0_t971 = 32'b00000000000000000000000000110000;
    FSM_fft_64_stage_6_0_t972 = FSM_fft_64_stage_6_0_t971[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t973 = 32'b00000000000000000000000000010000;
    FSM_fft_64_stage_6_0_t974 = FSM_fft_64_stage_6_0_t973[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t975 = i_data_in_imag[FSM_fft_64_stage_6_0_t974 * 32 +: 32];
    FSM_fft_64_stage_6_0_t976 = 32'b00000000000000000000000000110000;
    FSM_fft_64_stage_6_0_t977 = FSM_fft_64_stage_6_0_t976[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t978 = i_data_in_imag[FSM_fft_64_stage_6_0_t977 * 32 +: 32];
    FSM_fft_64_stage_6_0_t979 = FSM_fft_64_stage_6_0_t970;
    FSM_fft_64_stage_6_0_t979[FSM_fft_64_stage_6_0_t972 * 32 +: 32] = FSM_fft_64_stage_6_0_t975 - FSM_fft_64_stage_6_0_t978;
    FSM_fft_64_stage_6_0_t980 = 32'b00000000000000000000000000010001;
    FSM_fft_64_stage_6_0_t981 = FSM_fft_64_stage_6_0_t980[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t982 = 32'b00000000000000000000000000010001;
    FSM_fft_64_stage_6_0_t983 = FSM_fft_64_stage_6_0_t982[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t984 = i_data_in_imag[FSM_fft_64_stage_6_0_t983 * 32 +: 32];
    FSM_fft_64_stage_6_0_t985 = 32'b00000000000000000000000000110001;
    FSM_fft_64_stage_6_0_t986 = FSM_fft_64_stage_6_0_t985[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t987 = i_data_in_imag[FSM_fft_64_stage_6_0_t986 * 32 +: 32];
    FSM_fft_64_stage_6_0_t988 = FSM_fft_64_stage_6_0_t984 + FSM_fft_64_stage_6_0_t987;
    FSM_fft_64_stage_6_0_t989 = FSM_fft_64_stage_6_0_t988[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t990 = FSM_fft_64_stage_6_0_t979;
    FSM_fft_64_stage_6_0_t990[FSM_fft_64_stage_6_0_t981 * 32 +: 32] = FSM_fft_64_stage_6_0_t989;
    FSM_fft_64_stage_6_0_t991 = 32'b00000000000000000000000000110001;
    FSM_fft_64_stage_6_0_t992 = FSM_fft_64_stage_6_0_t991[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t993 = 32'b00000000000000000000000000010001;
    FSM_fft_64_stage_6_0_t994 = FSM_fft_64_stage_6_0_t993[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t995 = i_data_in_imag[FSM_fft_64_stage_6_0_t994 * 32 +: 32];
    FSM_fft_64_stage_6_0_t996 = 32'b00000000000000000000000000110001;
    FSM_fft_64_stage_6_0_t997 = FSM_fft_64_stage_6_0_t996[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t998 = i_data_in_imag[FSM_fft_64_stage_6_0_t997 * 32 +: 32];
    FSM_fft_64_stage_6_0_t999 = FSM_fft_64_stage_6_0_t990;
    FSM_fft_64_stage_6_0_t999[FSM_fft_64_stage_6_0_t992 * 32 +: 32] = FSM_fft_64_stage_6_0_t995 - FSM_fft_64_stage_6_0_t998;
    FSM_fft_64_stage_6_0_t1000 = 32'b00000000000000000000000000010010;
    FSM_fft_64_stage_6_0_t1001 = FSM_fft_64_stage_6_0_t1000[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1002 = 32'b00000000000000000000000000010010;
    FSM_fft_64_stage_6_0_t1003 = FSM_fft_64_stage_6_0_t1002[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1004 = i_data_in_imag[FSM_fft_64_stage_6_0_t1003 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1005 = 32'b00000000000000000000000000110010;
    FSM_fft_64_stage_6_0_t1006 = FSM_fft_64_stage_6_0_t1005[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1007 = i_data_in_imag[FSM_fft_64_stage_6_0_t1006 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1008 = FSM_fft_64_stage_6_0_t1004 + FSM_fft_64_stage_6_0_t1007;
    FSM_fft_64_stage_6_0_t1009 = FSM_fft_64_stage_6_0_t1008[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t1010 = FSM_fft_64_stage_6_0_t999;
    FSM_fft_64_stage_6_0_t1010[FSM_fft_64_stage_6_0_t1001 * 32 +: 32] = FSM_fft_64_stage_6_0_t1009;
    FSM_fft_64_stage_6_0_t1011 = 32'b00000000000000000000000000110010;
    FSM_fft_64_stage_6_0_t1012 = FSM_fft_64_stage_6_0_t1011[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1013 = 32'b00000000000000000000000000010010;
    FSM_fft_64_stage_6_0_t1014 = FSM_fft_64_stage_6_0_t1013[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1015 = i_data_in_imag[FSM_fft_64_stage_6_0_t1014 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1016 = 32'b00000000000000000000000000110010;
    FSM_fft_64_stage_6_0_t1017 = FSM_fft_64_stage_6_0_t1016[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1018 = i_data_in_imag[FSM_fft_64_stage_6_0_t1017 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1019 = FSM_fft_64_stage_6_0_t1010;
    FSM_fft_64_stage_6_0_t1019[FSM_fft_64_stage_6_0_t1012 * 32 +: 32] = FSM_fft_64_stage_6_0_t1015 - FSM_fft_64_stage_6_0_t1018;
    FSM_fft_64_stage_6_0_t1020 = 32'b00000000000000000000000000010011;
    FSM_fft_64_stage_6_0_t1021 = FSM_fft_64_stage_6_0_t1020[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1022 = 32'b00000000000000000000000000010011;
    FSM_fft_64_stage_6_0_t1023 = FSM_fft_64_stage_6_0_t1022[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1024 = i_data_in_imag[FSM_fft_64_stage_6_0_t1023 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1025 = 32'b00000000000000000000000000110011;
    FSM_fft_64_stage_6_0_t1026 = FSM_fft_64_stage_6_0_t1025[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1027 = i_data_in_imag[FSM_fft_64_stage_6_0_t1026 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1028 = FSM_fft_64_stage_6_0_t1024 + FSM_fft_64_stage_6_0_t1027;
    FSM_fft_64_stage_6_0_t1029 = FSM_fft_64_stage_6_0_t1028[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t1030 = FSM_fft_64_stage_6_0_t1019;
    FSM_fft_64_stage_6_0_t1030[FSM_fft_64_stage_6_0_t1021 * 32 +: 32] = FSM_fft_64_stage_6_0_t1029;
    FSM_fft_64_stage_6_0_t1031 = 32'b00000000000000000000000000110011;
    FSM_fft_64_stage_6_0_t1032 = FSM_fft_64_stage_6_0_t1031[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1033 = 32'b00000000000000000000000000010011;
    FSM_fft_64_stage_6_0_t1034 = FSM_fft_64_stage_6_0_t1033[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1035 = i_data_in_imag[FSM_fft_64_stage_6_0_t1034 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1036 = 32'b00000000000000000000000000110011;
    FSM_fft_64_stage_6_0_t1037 = FSM_fft_64_stage_6_0_t1036[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1038 = i_data_in_imag[FSM_fft_64_stage_6_0_t1037 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1039 = FSM_fft_64_stage_6_0_t1030;
    FSM_fft_64_stage_6_0_t1039[FSM_fft_64_stage_6_0_t1032 * 32 +: 32] = FSM_fft_64_stage_6_0_t1035 - FSM_fft_64_stage_6_0_t1038;
    FSM_fft_64_stage_6_0_t1040 = 32'b00000000000000000000000000010100;
    FSM_fft_64_stage_6_0_t1041 = FSM_fft_64_stage_6_0_t1040[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1042 = 32'b00000000000000000000000000010100;
    FSM_fft_64_stage_6_0_t1043 = FSM_fft_64_stage_6_0_t1042[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1044 = i_data_in_imag[FSM_fft_64_stage_6_0_t1043 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1045 = 32'b00000000000000000000000000110100;
    FSM_fft_64_stage_6_0_t1046 = FSM_fft_64_stage_6_0_t1045[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1047 = i_data_in_imag[FSM_fft_64_stage_6_0_t1046 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1048 = FSM_fft_64_stage_6_0_t1044 + FSM_fft_64_stage_6_0_t1047;
    FSM_fft_64_stage_6_0_t1049 = FSM_fft_64_stage_6_0_t1048[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t1050 = FSM_fft_64_stage_6_0_t1039;
    FSM_fft_64_stage_6_0_t1050[FSM_fft_64_stage_6_0_t1041 * 32 +: 32] = FSM_fft_64_stage_6_0_t1049;
    FSM_fft_64_stage_6_0_t1051 = 32'b00000000000000000000000000110100;
    FSM_fft_64_stage_6_0_t1052 = FSM_fft_64_stage_6_0_t1051[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1053 = 32'b00000000000000000000000000010100;
    FSM_fft_64_stage_6_0_t1054 = FSM_fft_64_stage_6_0_t1053[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1055 = i_data_in_imag[FSM_fft_64_stage_6_0_t1054 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1056 = 32'b00000000000000000000000000110100;
    FSM_fft_64_stage_6_0_t1057 = FSM_fft_64_stage_6_0_t1056[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1058 = i_data_in_imag[FSM_fft_64_stage_6_0_t1057 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1059 = FSM_fft_64_stage_6_0_t1050;
    FSM_fft_64_stage_6_0_t1059[FSM_fft_64_stage_6_0_t1052 * 32 +: 32] = FSM_fft_64_stage_6_0_t1055 - FSM_fft_64_stage_6_0_t1058;
    FSM_fft_64_stage_6_0_t1060 = 32'b00000000000000000000000000010101;
    FSM_fft_64_stage_6_0_t1061 = FSM_fft_64_stage_6_0_t1060[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1062 = 32'b00000000000000000000000000010101;
    FSM_fft_64_stage_6_0_t1063 = FSM_fft_64_stage_6_0_t1062[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1064 = i_data_in_imag[FSM_fft_64_stage_6_0_t1063 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1065 = 32'b00000000000000000000000000110101;
    FSM_fft_64_stage_6_0_t1066 = FSM_fft_64_stage_6_0_t1065[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1067 = i_data_in_imag[FSM_fft_64_stage_6_0_t1066 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1068 = FSM_fft_64_stage_6_0_t1064 + FSM_fft_64_stage_6_0_t1067;
    FSM_fft_64_stage_6_0_t1069 = FSM_fft_64_stage_6_0_t1068[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t1070 = FSM_fft_64_stage_6_0_t1059;
    FSM_fft_64_stage_6_0_t1070[FSM_fft_64_stage_6_0_t1061 * 32 +: 32] = FSM_fft_64_stage_6_0_t1069;
    FSM_fft_64_stage_6_0_t1071 = 32'b00000000000000000000000000110101;
    FSM_fft_64_stage_6_0_t1072 = FSM_fft_64_stage_6_0_t1071[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1073 = 32'b00000000000000000000000000010101;
    FSM_fft_64_stage_6_0_t1074 = FSM_fft_64_stage_6_0_t1073[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1075 = i_data_in_imag[FSM_fft_64_stage_6_0_t1074 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1076 = 32'b00000000000000000000000000110101;
    FSM_fft_64_stage_6_0_t1077 = FSM_fft_64_stage_6_0_t1076[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1078 = i_data_in_imag[FSM_fft_64_stage_6_0_t1077 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1079 = FSM_fft_64_stage_6_0_t1070;
    FSM_fft_64_stage_6_0_t1079[FSM_fft_64_stage_6_0_t1072 * 32 +: 32] = FSM_fft_64_stage_6_0_t1075 - FSM_fft_64_stage_6_0_t1078;
    FSM_fft_64_stage_6_0_t1080 = 32'b00000000000000000000000000010110;
    FSM_fft_64_stage_6_0_t1081 = FSM_fft_64_stage_6_0_t1080[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1082 = 32'b00000000000000000000000000010110;
    FSM_fft_64_stage_6_0_t1083 = FSM_fft_64_stage_6_0_t1082[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1084 = i_data_in_imag[FSM_fft_64_stage_6_0_t1083 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1085 = 32'b00000000000000000000000000110110;
    FSM_fft_64_stage_6_0_t1086 = FSM_fft_64_stage_6_0_t1085[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1087 = i_data_in_imag[FSM_fft_64_stage_6_0_t1086 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1088 = FSM_fft_64_stage_6_0_t1084 + FSM_fft_64_stage_6_0_t1087;
    FSM_fft_64_stage_6_0_t1089 = FSM_fft_64_stage_6_0_t1088[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t1090 = FSM_fft_64_stage_6_0_t1079;
    FSM_fft_64_stage_6_0_t1090[FSM_fft_64_stage_6_0_t1081 * 32 +: 32] = FSM_fft_64_stage_6_0_t1089;
    FSM_fft_64_stage_6_0_t1091 = 32'b00000000000000000000000000110110;
    FSM_fft_64_stage_6_0_t1092 = FSM_fft_64_stage_6_0_t1091[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1093 = 32'b00000000000000000000000000010110;
    FSM_fft_64_stage_6_0_t1094 = FSM_fft_64_stage_6_0_t1093[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1095 = i_data_in_imag[FSM_fft_64_stage_6_0_t1094 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1096 = 32'b00000000000000000000000000110110;
    FSM_fft_64_stage_6_0_t1097 = FSM_fft_64_stage_6_0_t1096[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1098 = i_data_in_imag[FSM_fft_64_stage_6_0_t1097 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1099 = FSM_fft_64_stage_6_0_t1090;
    FSM_fft_64_stage_6_0_t1099[FSM_fft_64_stage_6_0_t1092 * 32 +: 32] = FSM_fft_64_stage_6_0_t1095 - FSM_fft_64_stage_6_0_t1098;
    FSM_fft_64_stage_6_0_t1100 = 32'b00000000000000000000000000010111;
    FSM_fft_64_stage_6_0_t1101 = FSM_fft_64_stage_6_0_t1100[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1102 = 32'b00000000000000000000000000010111;
    FSM_fft_64_stage_6_0_t1103 = FSM_fft_64_stage_6_0_t1102[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1104 = i_data_in_imag[FSM_fft_64_stage_6_0_t1103 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1105 = 32'b00000000000000000000000000110111;
    FSM_fft_64_stage_6_0_t1106 = FSM_fft_64_stage_6_0_t1105[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1107 = i_data_in_imag[FSM_fft_64_stage_6_0_t1106 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1108 = FSM_fft_64_stage_6_0_t1104 + FSM_fft_64_stage_6_0_t1107;
    FSM_fft_64_stage_6_0_t1109 = FSM_fft_64_stage_6_0_t1108[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t1110 = FSM_fft_64_stage_6_0_t1099;
    FSM_fft_64_stage_6_0_t1110[FSM_fft_64_stage_6_0_t1101 * 32 +: 32] = FSM_fft_64_stage_6_0_t1109;
    FSM_fft_64_stage_6_0_t1111 = 32'b00000000000000000000000000110111;
    FSM_fft_64_stage_6_0_t1112 = FSM_fft_64_stage_6_0_t1111[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1113 = 32'b00000000000000000000000000010111;
    FSM_fft_64_stage_6_0_t1114 = FSM_fft_64_stage_6_0_t1113[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1115 = i_data_in_imag[FSM_fft_64_stage_6_0_t1114 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1116 = 32'b00000000000000000000000000110111;
    FSM_fft_64_stage_6_0_t1117 = FSM_fft_64_stage_6_0_t1116[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1118 = i_data_in_imag[FSM_fft_64_stage_6_0_t1117 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1119 = FSM_fft_64_stage_6_0_t1110;
    FSM_fft_64_stage_6_0_t1119[FSM_fft_64_stage_6_0_t1112 * 32 +: 32] = FSM_fft_64_stage_6_0_t1115 - FSM_fft_64_stage_6_0_t1118;
    FSM_fft_64_stage_6_0_t1120 = 32'b00000000000000000000000000011000;
    FSM_fft_64_stage_6_0_t1121 = FSM_fft_64_stage_6_0_t1120[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1122 = 32'b00000000000000000000000000011000;
    FSM_fft_64_stage_6_0_t1123 = FSM_fft_64_stage_6_0_t1122[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1124 = i_data_in_imag[FSM_fft_64_stage_6_0_t1123 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1125 = 32'b00000000000000000000000000111000;
    FSM_fft_64_stage_6_0_t1126 = FSM_fft_64_stage_6_0_t1125[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1127 = i_data_in_imag[FSM_fft_64_stage_6_0_t1126 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1128 = FSM_fft_64_stage_6_0_t1124 + FSM_fft_64_stage_6_0_t1127;
    FSM_fft_64_stage_6_0_t1129 = FSM_fft_64_stage_6_0_t1128[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t1130 = FSM_fft_64_stage_6_0_t1119;
    FSM_fft_64_stage_6_0_t1130[FSM_fft_64_stage_6_0_t1121 * 32 +: 32] = FSM_fft_64_stage_6_0_t1129;
    FSM_fft_64_stage_6_0_t1131 = 32'b00000000000000000000000000111000;
    FSM_fft_64_stage_6_0_t1132 = FSM_fft_64_stage_6_0_t1131[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1133 = 32'b00000000000000000000000000011000;
    FSM_fft_64_stage_6_0_t1134 = FSM_fft_64_stage_6_0_t1133[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1135 = i_data_in_imag[FSM_fft_64_stage_6_0_t1134 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1136 = 32'b00000000000000000000000000111000;
    FSM_fft_64_stage_6_0_t1137 = FSM_fft_64_stage_6_0_t1136[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1138 = i_data_in_imag[FSM_fft_64_stage_6_0_t1137 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1139 = FSM_fft_64_stage_6_0_t1130;
    FSM_fft_64_stage_6_0_t1139[FSM_fft_64_stage_6_0_t1132 * 32 +: 32] = FSM_fft_64_stage_6_0_t1135 - FSM_fft_64_stage_6_0_t1138;
    FSM_fft_64_stage_6_0_t1140 = 32'b00000000000000000000000000011001;
    FSM_fft_64_stage_6_0_t1141 = FSM_fft_64_stage_6_0_t1140[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1142 = 32'b00000000000000000000000000011001;
    FSM_fft_64_stage_6_0_t1143 = FSM_fft_64_stage_6_0_t1142[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1144 = i_data_in_imag[FSM_fft_64_stage_6_0_t1143 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1145 = 32'b00000000000000000000000000111001;
    FSM_fft_64_stage_6_0_t1146 = FSM_fft_64_stage_6_0_t1145[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1147 = i_data_in_imag[FSM_fft_64_stage_6_0_t1146 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1148 = FSM_fft_64_stage_6_0_t1144 + FSM_fft_64_stage_6_0_t1147;
    FSM_fft_64_stage_6_0_t1149 = FSM_fft_64_stage_6_0_t1148[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t1150 = FSM_fft_64_stage_6_0_t1139;
    FSM_fft_64_stage_6_0_t1150[FSM_fft_64_stage_6_0_t1141 * 32 +: 32] = FSM_fft_64_stage_6_0_t1149;
    FSM_fft_64_stage_6_0_t1151 = 32'b00000000000000000000000000111001;
    FSM_fft_64_stage_6_0_t1152 = FSM_fft_64_stage_6_0_t1151[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1153 = 32'b00000000000000000000000000011001;
    FSM_fft_64_stage_6_0_t1154 = FSM_fft_64_stage_6_0_t1153[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1155 = i_data_in_imag[FSM_fft_64_stage_6_0_t1154 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1156 = 32'b00000000000000000000000000111001;
    FSM_fft_64_stage_6_0_t1157 = FSM_fft_64_stage_6_0_t1156[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1158 = i_data_in_imag[FSM_fft_64_stage_6_0_t1157 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1159 = FSM_fft_64_stage_6_0_t1150;
    FSM_fft_64_stage_6_0_t1159[FSM_fft_64_stage_6_0_t1152 * 32 +: 32] = FSM_fft_64_stage_6_0_t1155 - FSM_fft_64_stage_6_0_t1158;
    FSM_fft_64_stage_6_0_t1160 = 32'b00000000000000000000000000011010;
    FSM_fft_64_stage_6_0_t1161 = FSM_fft_64_stage_6_0_t1160[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1162 = 32'b00000000000000000000000000011010;
    FSM_fft_64_stage_6_0_t1163 = FSM_fft_64_stage_6_0_t1162[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1164 = i_data_in_imag[FSM_fft_64_stage_6_0_t1163 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1165 = 32'b00000000000000000000000000111010;
    FSM_fft_64_stage_6_0_t1166 = FSM_fft_64_stage_6_0_t1165[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1167 = i_data_in_imag[FSM_fft_64_stage_6_0_t1166 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1168 = FSM_fft_64_stage_6_0_t1164 + FSM_fft_64_stage_6_0_t1167;
    FSM_fft_64_stage_6_0_t1169 = FSM_fft_64_stage_6_0_t1168[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t1170 = FSM_fft_64_stage_6_0_t1159;
    FSM_fft_64_stage_6_0_t1170[FSM_fft_64_stage_6_0_t1161 * 32 +: 32] = FSM_fft_64_stage_6_0_t1169;
    FSM_fft_64_stage_6_0_t1171 = 32'b00000000000000000000000000111010;
    FSM_fft_64_stage_6_0_t1172 = FSM_fft_64_stage_6_0_t1171[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1173 = 32'b00000000000000000000000000011010;
    FSM_fft_64_stage_6_0_t1174 = FSM_fft_64_stage_6_0_t1173[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1175 = i_data_in_imag[FSM_fft_64_stage_6_0_t1174 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1176 = 32'b00000000000000000000000000111010;
    FSM_fft_64_stage_6_0_t1177 = FSM_fft_64_stage_6_0_t1176[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1178 = i_data_in_imag[FSM_fft_64_stage_6_0_t1177 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1179 = FSM_fft_64_stage_6_0_t1170;
    FSM_fft_64_stage_6_0_t1179[FSM_fft_64_stage_6_0_t1172 * 32 +: 32] = FSM_fft_64_stage_6_0_t1175 - FSM_fft_64_stage_6_0_t1178;
    FSM_fft_64_stage_6_0_t1180 = 32'b00000000000000000000000000011011;
    FSM_fft_64_stage_6_0_t1181 = FSM_fft_64_stage_6_0_t1180[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1182 = 32'b00000000000000000000000000011011;
    FSM_fft_64_stage_6_0_t1183 = FSM_fft_64_stage_6_0_t1182[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1184 = i_data_in_imag[FSM_fft_64_stage_6_0_t1183 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1185 = 32'b00000000000000000000000000111011;
    FSM_fft_64_stage_6_0_t1186 = FSM_fft_64_stage_6_0_t1185[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1187 = i_data_in_imag[FSM_fft_64_stage_6_0_t1186 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1188 = FSM_fft_64_stage_6_0_t1184 + FSM_fft_64_stage_6_0_t1187;
    FSM_fft_64_stage_6_0_t1189 = FSM_fft_64_stage_6_0_t1188[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t1190 = FSM_fft_64_stage_6_0_t1179;
    FSM_fft_64_stage_6_0_t1190[FSM_fft_64_stage_6_0_t1181 * 32 +: 32] = FSM_fft_64_stage_6_0_t1189;
    FSM_fft_64_stage_6_0_t1191 = 32'b00000000000000000000000000111011;
    FSM_fft_64_stage_6_0_t1192 = FSM_fft_64_stage_6_0_t1191[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1193 = 32'b00000000000000000000000000011011;
    FSM_fft_64_stage_6_0_t1194 = FSM_fft_64_stage_6_0_t1193[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1195 = i_data_in_imag[FSM_fft_64_stage_6_0_t1194 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1196 = 32'b00000000000000000000000000111011;
    FSM_fft_64_stage_6_0_t1197 = FSM_fft_64_stage_6_0_t1196[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1198 = i_data_in_imag[FSM_fft_64_stage_6_0_t1197 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1199 = FSM_fft_64_stage_6_0_t1190;
    FSM_fft_64_stage_6_0_t1199[FSM_fft_64_stage_6_0_t1192 * 32 +: 32] = FSM_fft_64_stage_6_0_t1195 - FSM_fft_64_stage_6_0_t1198;
    FSM_fft_64_stage_6_0_t1200 = 32'b00000000000000000000000000011100;
    FSM_fft_64_stage_6_0_t1201 = FSM_fft_64_stage_6_0_t1200[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1202 = 32'b00000000000000000000000000011100;
    FSM_fft_64_stage_6_0_t1203 = FSM_fft_64_stage_6_0_t1202[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1204 = i_data_in_imag[FSM_fft_64_stage_6_0_t1203 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1205 = 32'b00000000000000000000000000111100;
    FSM_fft_64_stage_6_0_t1206 = FSM_fft_64_stage_6_0_t1205[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1207 = i_data_in_imag[FSM_fft_64_stage_6_0_t1206 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1208 = FSM_fft_64_stage_6_0_t1204 + FSM_fft_64_stage_6_0_t1207;
    FSM_fft_64_stage_6_0_t1209 = FSM_fft_64_stage_6_0_t1208[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t1210 = FSM_fft_64_stage_6_0_t1199;
    FSM_fft_64_stage_6_0_t1210[FSM_fft_64_stage_6_0_t1201 * 32 +: 32] = FSM_fft_64_stage_6_0_t1209;
    FSM_fft_64_stage_6_0_t1211 = 32'b00000000000000000000000000111100;
    FSM_fft_64_stage_6_0_t1212 = FSM_fft_64_stage_6_0_t1211[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1213 = 32'b00000000000000000000000000011100;
    FSM_fft_64_stage_6_0_t1214 = FSM_fft_64_stage_6_0_t1213[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1215 = i_data_in_imag[FSM_fft_64_stage_6_0_t1214 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1216 = 32'b00000000000000000000000000111100;
    FSM_fft_64_stage_6_0_t1217 = FSM_fft_64_stage_6_0_t1216[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1218 = i_data_in_imag[FSM_fft_64_stage_6_0_t1217 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1219 = FSM_fft_64_stage_6_0_t1210;
    FSM_fft_64_stage_6_0_t1219[FSM_fft_64_stage_6_0_t1212 * 32 +: 32] = FSM_fft_64_stage_6_0_t1215 - FSM_fft_64_stage_6_0_t1218;
    FSM_fft_64_stage_6_0_t1220 = 32'b00000000000000000000000000011101;
    FSM_fft_64_stage_6_0_t1221 = FSM_fft_64_stage_6_0_t1220[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1222 = 32'b00000000000000000000000000011101;
    FSM_fft_64_stage_6_0_t1223 = FSM_fft_64_stage_6_0_t1222[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1224 = i_data_in_imag[FSM_fft_64_stage_6_0_t1223 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1225 = 32'b00000000000000000000000000111101;
    FSM_fft_64_stage_6_0_t1226 = FSM_fft_64_stage_6_0_t1225[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1227 = i_data_in_imag[FSM_fft_64_stage_6_0_t1226 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1228 = FSM_fft_64_stage_6_0_t1224 + FSM_fft_64_stage_6_0_t1227;
    FSM_fft_64_stage_6_0_t1229 = FSM_fft_64_stage_6_0_t1228[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t1230 = FSM_fft_64_stage_6_0_t1219;
    FSM_fft_64_stage_6_0_t1230[FSM_fft_64_stage_6_0_t1221 * 32 +: 32] = FSM_fft_64_stage_6_0_t1229;
    FSM_fft_64_stage_6_0_t1231 = 32'b00000000000000000000000000111101;
    FSM_fft_64_stage_6_0_t1232 = FSM_fft_64_stage_6_0_t1231[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1233 = 32'b00000000000000000000000000011101;
    FSM_fft_64_stage_6_0_t1234 = FSM_fft_64_stage_6_0_t1233[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1235 = i_data_in_imag[FSM_fft_64_stage_6_0_t1234 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1236 = 32'b00000000000000000000000000111101;
    FSM_fft_64_stage_6_0_t1237 = FSM_fft_64_stage_6_0_t1236[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1238 = i_data_in_imag[FSM_fft_64_stage_6_0_t1237 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1239 = FSM_fft_64_stage_6_0_t1230;
    FSM_fft_64_stage_6_0_t1239[FSM_fft_64_stage_6_0_t1232 * 32 +: 32] = FSM_fft_64_stage_6_0_t1235 - FSM_fft_64_stage_6_0_t1238;
    FSM_fft_64_stage_6_0_t1240 = 32'b00000000000000000000000000011110;
    FSM_fft_64_stage_6_0_t1241 = FSM_fft_64_stage_6_0_t1240[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1242 = 32'b00000000000000000000000000011110;
    FSM_fft_64_stage_6_0_t1243 = FSM_fft_64_stage_6_0_t1242[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1244 = i_data_in_imag[FSM_fft_64_stage_6_0_t1243 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1245 = 32'b00000000000000000000000000111110;
    FSM_fft_64_stage_6_0_t1246 = FSM_fft_64_stage_6_0_t1245[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1247 = i_data_in_imag[FSM_fft_64_stage_6_0_t1246 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1248 = FSM_fft_64_stage_6_0_t1244 + FSM_fft_64_stage_6_0_t1247;
    FSM_fft_64_stage_6_0_t1249 = FSM_fft_64_stage_6_0_t1248[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t1250 = FSM_fft_64_stage_6_0_t1239;
    FSM_fft_64_stage_6_0_t1250[FSM_fft_64_stage_6_0_t1241 * 32 +: 32] = FSM_fft_64_stage_6_0_t1249;
    FSM_fft_64_stage_6_0_t1251 = 32'b00000000000000000000000000111110;
    FSM_fft_64_stage_6_0_t1252 = FSM_fft_64_stage_6_0_t1251[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1253 = 32'b00000000000000000000000000011110;
    FSM_fft_64_stage_6_0_t1254 = FSM_fft_64_stage_6_0_t1253[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1255 = i_data_in_imag[FSM_fft_64_stage_6_0_t1254 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1256 = 32'b00000000000000000000000000111110;
    FSM_fft_64_stage_6_0_t1257 = FSM_fft_64_stage_6_0_t1256[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1258 = i_data_in_imag[FSM_fft_64_stage_6_0_t1257 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1259 = FSM_fft_64_stage_6_0_t1250;
    FSM_fft_64_stage_6_0_t1259[FSM_fft_64_stage_6_0_t1252 * 32 +: 32] = FSM_fft_64_stage_6_0_t1255 - FSM_fft_64_stage_6_0_t1258;
    FSM_fft_64_stage_6_0_t1260 = 32'b00000000000000000000000000011111;
    FSM_fft_64_stage_6_0_t1261 = FSM_fft_64_stage_6_0_t1260[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1262 = 32'b00000000000000000000000000011111;
    FSM_fft_64_stage_6_0_t1263 = FSM_fft_64_stage_6_0_t1262[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1264 = i_data_in_imag[FSM_fft_64_stage_6_0_t1263 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1265 = 32'b00000000000000000000000000111111;
    FSM_fft_64_stage_6_0_t1266 = FSM_fft_64_stage_6_0_t1265[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1267 = i_data_in_imag[FSM_fft_64_stage_6_0_t1266 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1268 = FSM_fft_64_stage_6_0_t1264 + FSM_fft_64_stage_6_0_t1267;
    FSM_fft_64_stage_6_0_t1269 = FSM_fft_64_stage_6_0_t1268[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t1270 = FSM_fft_64_stage_6_0_t1259;
    FSM_fft_64_stage_6_0_t1270[FSM_fft_64_stage_6_0_t1261 * 32 +: 32] = FSM_fft_64_stage_6_0_t1269;
    FSM_fft_64_stage_6_0_t1271 = 32'b00000000000000000000000000111111;
    FSM_fft_64_stage_6_0_t1272 = FSM_fft_64_stage_6_0_t1271[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1273 = 32'b00000000000000000000000000011111;
    FSM_fft_64_stage_6_0_t1274 = FSM_fft_64_stage_6_0_t1273[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1275 = i_data_in_imag[FSM_fft_64_stage_6_0_t1274 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1276 = 32'b00000000000000000000000000111111;
    FSM_fft_64_stage_6_0_t1277 = FSM_fft_64_stage_6_0_t1276[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1278 = i_data_in_imag[FSM_fft_64_stage_6_0_t1277 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1279 = FSM_fft_64_stage_6_0_t1270;
    FSM_fft_64_stage_6_0_t1279[FSM_fft_64_stage_6_0_t1272 * 32 +: 32] = FSM_fft_64_stage_6_0_t1275 - FSM_fft_64_stage_6_0_t1278;
end

always @* begin
    FSM_fft_64_stage_6_0_t0 = 32'b0;
    FSM_fft_64_stage_6_0_t1 = FSM_fft_64_stage_6_0_t0[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t2 = 32'b0;
    FSM_fft_64_stage_6_0_t3 = FSM_fft_64_stage_6_0_t2[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t4 = i_data_in_real[FSM_fft_64_stage_6_0_t3 * 32 +: 32];
    FSM_fft_64_stage_6_0_t5 = 32'b00000000000000000000000000100000;
    FSM_fft_64_stage_6_0_t6 = FSM_fft_64_stage_6_0_t5[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t7 = i_data_in_real[FSM_fft_64_stage_6_0_t6 * 32 +: 32];
    FSM_fft_64_stage_6_0_t8 = FSM_fft_64_stage_6_0_t4 + FSM_fft_64_stage_6_0_t7;
    FSM_fft_64_stage_6_0_t9 = FSM_fft_64_stage_6_0_t8[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t10 = i_data_in_real;
    FSM_fft_64_stage_6_0_t10[FSM_fft_64_stage_6_0_t1 * 32 +: 32] = FSM_fft_64_stage_6_0_t9;
    FSM_fft_64_stage_6_0_t11 = 32'b00000000000000000000000000100000;
    FSM_fft_64_stage_6_0_t12 = FSM_fft_64_stage_6_0_t11[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t13 = 32'b0;
    FSM_fft_64_stage_6_0_t14 = FSM_fft_64_stage_6_0_t13[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t15 = i_data_in_real[FSM_fft_64_stage_6_0_t14 * 32 +: 32];
    FSM_fft_64_stage_6_0_t16 = 32'b00000000000000000000000000100000;
    FSM_fft_64_stage_6_0_t17 = FSM_fft_64_stage_6_0_t16[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t18 = i_data_in_real[FSM_fft_64_stage_6_0_t17 * 32 +: 32];
    FSM_fft_64_stage_6_0_t19 = FSM_fft_64_stage_6_0_t10;
    FSM_fft_64_stage_6_0_t19[FSM_fft_64_stage_6_0_t12 * 32 +: 32] = FSM_fft_64_stage_6_0_t15 - FSM_fft_64_stage_6_0_t18;
    FSM_fft_64_stage_6_0_t20 = 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_6_0_t21 = FSM_fft_64_stage_6_0_t20[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t22 = 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_6_0_t23 = FSM_fft_64_stage_6_0_t22[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t24 = i_data_in_real[FSM_fft_64_stage_6_0_t23 * 32 +: 32];
    FSM_fft_64_stage_6_0_t25 = 32'b00000000000000000000000000100001;
    FSM_fft_64_stage_6_0_t26 = FSM_fft_64_stage_6_0_t25[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t27 = i_data_in_real[FSM_fft_64_stage_6_0_t26 * 32 +: 32];
    FSM_fft_64_stage_6_0_t28 = FSM_fft_64_stage_6_0_t24 + FSM_fft_64_stage_6_0_t27;
    FSM_fft_64_stage_6_0_t29 = FSM_fft_64_stage_6_0_t28[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t30 = FSM_fft_64_stage_6_0_t19;
    FSM_fft_64_stage_6_0_t30[FSM_fft_64_stage_6_0_t21 * 32 +: 32] = FSM_fft_64_stage_6_0_t29;
    FSM_fft_64_stage_6_0_t31 = 32'b00000000000000000000000000100001;
    FSM_fft_64_stage_6_0_t32 = FSM_fft_64_stage_6_0_t31[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t33 = 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_6_0_t34 = FSM_fft_64_stage_6_0_t33[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t35 = i_data_in_real[FSM_fft_64_stage_6_0_t34 * 32 +: 32];
    FSM_fft_64_stage_6_0_t36 = 32'b00000000000000000000000000100001;
    FSM_fft_64_stage_6_0_t37 = FSM_fft_64_stage_6_0_t36[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t38 = i_data_in_real[FSM_fft_64_stage_6_0_t37 * 32 +: 32];
    FSM_fft_64_stage_6_0_t39 = FSM_fft_64_stage_6_0_t30;
    FSM_fft_64_stage_6_0_t39[FSM_fft_64_stage_6_0_t32 * 32 +: 32] = FSM_fft_64_stage_6_0_t35 - FSM_fft_64_stage_6_0_t38;
    FSM_fft_64_stage_6_0_t40 = 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_6_0_t41 = FSM_fft_64_stage_6_0_t40[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t42 = 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_6_0_t43 = FSM_fft_64_stage_6_0_t42[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t44 = i_data_in_real[FSM_fft_64_stage_6_0_t43 * 32 +: 32];
    FSM_fft_64_stage_6_0_t45 = 32'b00000000000000000000000000100010;
    FSM_fft_64_stage_6_0_t46 = FSM_fft_64_stage_6_0_t45[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t47 = i_data_in_real[FSM_fft_64_stage_6_0_t46 * 32 +: 32];
    FSM_fft_64_stage_6_0_t48 = FSM_fft_64_stage_6_0_t44 + FSM_fft_64_stage_6_0_t47;
    FSM_fft_64_stage_6_0_t49 = FSM_fft_64_stage_6_0_t48[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t50 = FSM_fft_64_stage_6_0_t39;
    FSM_fft_64_stage_6_0_t50[FSM_fft_64_stage_6_0_t41 * 32 +: 32] = FSM_fft_64_stage_6_0_t49;
    FSM_fft_64_stage_6_0_t51 = 32'b00000000000000000000000000100010;
    FSM_fft_64_stage_6_0_t52 = FSM_fft_64_stage_6_0_t51[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t53 = 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_6_0_t54 = FSM_fft_64_stage_6_0_t53[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t55 = i_data_in_real[FSM_fft_64_stage_6_0_t54 * 32 +: 32];
    FSM_fft_64_stage_6_0_t56 = 32'b00000000000000000000000000100010;
    FSM_fft_64_stage_6_0_t57 = FSM_fft_64_stage_6_0_t56[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t58 = i_data_in_real[FSM_fft_64_stage_6_0_t57 * 32 +: 32];
    FSM_fft_64_stage_6_0_t59 = FSM_fft_64_stage_6_0_t50;
    FSM_fft_64_stage_6_0_t59[FSM_fft_64_stage_6_0_t52 * 32 +: 32] = FSM_fft_64_stage_6_0_t55 - FSM_fft_64_stage_6_0_t58;
    FSM_fft_64_stage_6_0_t60 = 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_6_0_t61 = FSM_fft_64_stage_6_0_t60[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t62 = 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_6_0_t63 = FSM_fft_64_stage_6_0_t62[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t64 = i_data_in_real[FSM_fft_64_stage_6_0_t63 * 32 +: 32];
    FSM_fft_64_stage_6_0_t65 = 32'b00000000000000000000000000100011;
    FSM_fft_64_stage_6_0_t66 = FSM_fft_64_stage_6_0_t65[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t67 = i_data_in_real[FSM_fft_64_stage_6_0_t66 * 32 +: 32];
    FSM_fft_64_stage_6_0_t68 = FSM_fft_64_stage_6_0_t64 + FSM_fft_64_stage_6_0_t67;
    FSM_fft_64_stage_6_0_t69 = FSM_fft_64_stage_6_0_t68[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t70 = FSM_fft_64_stage_6_0_t59;
    FSM_fft_64_stage_6_0_t70[FSM_fft_64_stage_6_0_t61 * 32 +: 32] = FSM_fft_64_stage_6_0_t69;
    FSM_fft_64_stage_6_0_t71 = 32'b00000000000000000000000000100011;
    FSM_fft_64_stage_6_0_t72 = FSM_fft_64_stage_6_0_t71[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t73 = 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_6_0_t74 = FSM_fft_64_stage_6_0_t73[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t75 = i_data_in_real[FSM_fft_64_stage_6_0_t74 * 32 +: 32];
    FSM_fft_64_stage_6_0_t76 = 32'b00000000000000000000000000100011;
    FSM_fft_64_stage_6_0_t77 = FSM_fft_64_stage_6_0_t76[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t78 = i_data_in_real[FSM_fft_64_stage_6_0_t77 * 32 +: 32];
    FSM_fft_64_stage_6_0_t79 = FSM_fft_64_stage_6_0_t70;
    FSM_fft_64_stage_6_0_t79[FSM_fft_64_stage_6_0_t72 * 32 +: 32] = FSM_fft_64_stage_6_0_t75 - FSM_fft_64_stage_6_0_t78;
    FSM_fft_64_stage_6_0_t80 = 32'b00000000000000000000000000000100;
    FSM_fft_64_stage_6_0_t81 = FSM_fft_64_stage_6_0_t80[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t82 = 32'b00000000000000000000000000000100;
    FSM_fft_64_stage_6_0_t83 = FSM_fft_64_stage_6_0_t82[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t84 = i_data_in_real[FSM_fft_64_stage_6_0_t83 * 32 +: 32];
    FSM_fft_64_stage_6_0_t85 = 32'b00000000000000000000000000100100;
    FSM_fft_64_stage_6_0_t86 = FSM_fft_64_stage_6_0_t85[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t87 = i_data_in_real[FSM_fft_64_stage_6_0_t86 * 32 +: 32];
    FSM_fft_64_stage_6_0_t88 = FSM_fft_64_stage_6_0_t84 + FSM_fft_64_stage_6_0_t87;
    FSM_fft_64_stage_6_0_t89 = FSM_fft_64_stage_6_0_t88[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t90 = FSM_fft_64_stage_6_0_t79;
    FSM_fft_64_stage_6_0_t90[FSM_fft_64_stage_6_0_t81 * 32 +: 32] = FSM_fft_64_stage_6_0_t89;
    FSM_fft_64_stage_6_0_t91 = 32'b00000000000000000000000000100100;
    FSM_fft_64_stage_6_0_t92 = FSM_fft_64_stage_6_0_t91[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t93 = 32'b00000000000000000000000000000100;
    FSM_fft_64_stage_6_0_t94 = FSM_fft_64_stage_6_0_t93[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t95 = i_data_in_real[FSM_fft_64_stage_6_0_t94 * 32 +: 32];
    FSM_fft_64_stage_6_0_t96 = 32'b00000000000000000000000000100100;
    FSM_fft_64_stage_6_0_t97 = FSM_fft_64_stage_6_0_t96[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t98 = i_data_in_real[FSM_fft_64_stage_6_0_t97 * 32 +: 32];
    FSM_fft_64_stage_6_0_t99 = FSM_fft_64_stage_6_0_t90;
    FSM_fft_64_stage_6_0_t99[FSM_fft_64_stage_6_0_t92 * 32 +: 32] = FSM_fft_64_stage_6_0_t95 - FSM_fft_64_stage_6_0_t98;
    FSM_fft_64_stage_6_0_t100 = 32'b00000000000000000000000000000101;
    FSM_fft_64_stage_6_0_t101 = FSM_fft_64_stage_6_0_t100[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t102 = 32'b00000000000000000000000000000101;
    FSM_fft_64_stage_6_0_t103 = FSM_fft_64_stage_6_0_t102[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t104 = i_data_in_real[FSM_fft_64_stage_6_0_t103 * 32 +: 32];
    FSM_fft_64_stage_6_0_t105 = 32'b00000000000000000000000000100101;
    FSM_fft_64_stage_6_0_t106 = FSM_fft_64_stage_6_0_t105[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t107 = i_data_in_real[FSM_fft_64_stage_6_0_t106 * 32 +: 32];
    FSM_fft_64_stage_6_0_t108 = FSM_fft_64_stage_6_0_t104 + FSM_fft_64_stage_6_0_t107;
    FSM_fft_64_stage_6_0_t109 = FSM_fft_64_stage_6_0_t108[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t110 = FSM_fft_64_stage_6_0_t99;
    FSM_fft_64_stage_6_0_t110[FSM_fft_64_stage_6_0_t101 * 32 +: 32] = FSM_fft_64_stage_6_0_t109;
    FSM_fft_64_stage_6_0_t111 = 32'b00000000000000000000000000100101;
    FSM_fft_64_stage_6_0_t112 = FSM_fft_64_stage_6_0_t111[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t113 = 32'b00000000000000000000000000000101;
    FSM_fft_64_stage_6_0_t114 = FSM_fft_64_stage_6_0_t113[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t115 = i_data_in_real[FSM_fft_64_stage_6_0_t114 * 32 +: 32];
    FSM_fft_64_stage_6_0_t116 = 32'b00000000000000000000000000100101;
    FSM_fft_64_stage_6_0_t117 = FSM_fft_64_stage_6_0_t116[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t118 = i_data_in_real[FSM_fft_64_stage_6_0_t117 * 32 +: 32];
    FSM_fft_64_stage_6_0_t119 = FSM_fft_64_stage_6_0_t110;
    FSM_fft_64_stage_6_0_t119[FSM_fft_64_stage_6_0_t112 * 32 +: 32] = FSM_fft_64_stage_6_0_t115 - FSM_fft_64_stage_6_0_t118;
    FSM_fft_64_stage_6_0_t120 = 32'b00000000000000000000000000000110;
    FSM_fft_64_stage_6_0_t121 = FSM_fft_64_stage_6_0_t120[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t122 = 32'b00000000000000000000000000000110;
    FSM_fft_64_stage_6_0_t123 = FSM_fft_64_stage_6_0_t122[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t124 = i_data_in_real[FSM_fft_64_stage_6_0_t123 * 32 +: 32];
    FSM_fft_64_stage_6_0_t125 = 32'b00000000000000000000000000100110;
    FSM_fft_64_stage_6_0_t126 = FSM_fft_64_stage_6_0_t125[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t127 = i_data_in_real[FSM_fft_64_stage_6_0_t126 * 32 +: 32];
    FSM_fft_64_stage_6_0_t128 = FSM_fft_64_stage_6_0_t124 + FSM_fft_64_stage_6_0_t127;
    FSM_fft_64_stage_6_0_t129 = FSM_fft_64_stage_6_0_t128[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t130 = FSM_fft_64_stage_6_0_t119;
    FSM_fft_64_stage_6_0_t130[FSM_fft_64_stage_6_0_t121 * 32 +: 32] = FSM_fft_64_stage_6_0_t129;
    FSM_fft_64_stage_6_0_t131 = 32'b00000000000000000000000000100110;
    FSM_fft_64_stage_6_0_t132 = FSM_fft_64_stage_6_0_t131[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t133 = 32'b00000000000000000000000000000110;
    FSM_fft_64_stage_6_0_t134 = FSM_fft_64_stage_6_0_t133[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t135 = i_data_in_real[FSM_fft_64_stage_6_0_t134 * 32 +: 32];
    FSM_fft_64_stage_6_0_t136 = 32'b00000000000000000000000000100110;
    FSM_fft_64_stage_6_0_t137 = FSM_fft_64_stage_6_0_t136[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t138 = i_data_in_real[FSM_fft_64_stage_6_0_t137 * 32 +: 32];
    FSM_fft_64_stage_6_0_t139 = FSM_fft_64_stage_6_0_t130;
    FSM_fft_64_stage_6_0_t139[FSM_fft_64_stage_6_0_t132 * 32 +: 32] = FSM_fft_64_stage_6_0_t135 - FSM_fft_64_stage_6_0_t138;
    FSM_fft_64_stage_6_0_t140 = 32'b00000000000000000000000000000111;
    FSM_fft_64_stage_6_0_t141 = FSM_fft_64_stage_6_0_t140[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t142 = 32'b00000000000000000000000000000111;
    FSM_fft_64_stage_6_0_t143 = FSM_fft_64_stage_6_0_t142[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t144 = i_data_in_real[FSM_fft_64_stage_6_0_t143 * 32 +: 32];
    FSM_fft_64_stage_6_0_t145 = 32'b00000000000000000000000000100111;
    FSM_fft_64_stage_6_0_t146 = FSM_fft_64_stage_6_0_t145[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t147 = i_data_in_real[FSM_fft_64_stage_6_0_t146 * 32 +: 32];
    FSM_fft_64_stage_6_0_t148 = FSM_fft_64_stage_6_0_t144 + FSM_fft_64_stage_6_0_t147;
    FSM_fft_64_stage_6_0_t149 = FSM_fft_64_stage_6_0_t148[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t150 = FSM_fft_64_stage_6_0_t139;
    FSM_fft_64_stage_6_0_t150[FSM_fft_64_stage_6_0_t141 * 32 +: 32] = FSM_fft_64_stage_6_0_t149;
    FSM_fft_64_stage_6_0_t151 = 32'b00000000000000000000000000100111;
    FSM_fft_64_stage_6_0_t152 = FSM_fft_64_stage_6_0_t151[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t153 = 32'b00000000000000000000000000000111;
    FSM_fft_64_stage_6_0_t154 = FSM_fft_64_stage_6_0_t153[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t155 = i_data_in_real[FSM_fft_64_stage_6_0_t154 * 32 +: 32];
    FSM_fft_64_stage_6_0_t156 = 32'b00000000000000000000000000100111;
    FSM_fft_64_stage_6_0_t157 = FSM_fft_64_stage_6_0_t156[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t158 = i_data_in_real[FSM_fft_64_stage_6_0_t157 * 32 +: 32];
    FSM_fft_64_stage_6_0_t159 = FSM_fft_64_stage_6_0_t150;
    FSM_fft_64_stage_6_0_t159[FSM_fft_64_stage_6_0_t152 * 32 +: 32] = FSM_fft_64_stage_6_0_t155 - FSM_fft_64_stage_6_0_t158;
    FSM_fft_64_stage_6_0_t160 = 32'b00000000000000000000000000001000;
    FSM_fft_64_stage_6_0_t161 = FSM_fft_64_stage_6_0_t160[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t162 = 32'b00000000000000000000000000001000;
    FSM_fft_64_stage_6_0_t163 = FSM_fft_64_stage_6_0_t162[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t164 = i_data_in_real[FSM_fft_64_stage_6_0_t163 * 32 +: 32];
    FSM_fft_64_stage_6_0_t165 = 32'b00000000000000000000000000101000;
    FSM_fft_64_stage_6_0_t166 = FSM_fft_64_stage_6_0_t165[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t167 = i_data_in_real[FSM_fft_64_stage_6_0_t166 * 32 +: 32];
    FSM_fft_64_stage_6_0_t168 = FSM_fft_64_stage_6_0_t164 + FSM_fft_64_stage_6_0_t167;
    FSM_fft_64_stage_6_0_t169 = FSM_fft_64_stage_6_0_t168[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t170 = FSM_fft_64_stage_6_0_t159;
    FSM_fft_64_stage_6_0_t170[FSM_fft_64_stage_6_0_t161 * 32 +: 32] = FSM_fft_64_stage_6_0_t169;
    FSM_fft_64_stage_6_0_t171 = 32'b00000000000000000000000000101000;
    FSM_fft_64_stage_6_0_t172 = FSM_fft_64_stage_6_0_t171[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t173 = 32'b00000000000000000000000000001000;
    FSM_fft_64_stage_6_0_t174 = FSM_fft_64_stage_6_0_t173[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t175 = i_data_in_real[FSM_fft_64_stage_6_0_t174 * 32 +: 32];
    FSM_fft_64_stage_6_0_t176 = 32'b00000000000000000000000000101000;
    FSM_fft_64_stage_6_0_t177 = FSM_fft_64_stage_6_0_t176[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t178 = i_data_in_real[FSM_fft_64_stage_6_0_t177 * 32 +: 32];
    FSM_fft_64_stage_6_0_t179 = FSM_fft_64_stage_6_0_t170;
    FSM_fft_64_stage_6_0_t179[FSM_fft_64_stage_6_0_t172 * 32 +: 32] = FSM_fft_64_stage_6_0_t175 - FSM_fft_64_stage_6_0_t178;
    FSM_fft_64_stage_6_0_t180 = 32'b00000000000000000000000000001001;
    FSM_fft_64_stage_6_0_t181 = FSM_fft_64_stage_6_0_t180[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t182 = 32'b00000000000000000000000000001001;
    FSM_fft_64_stage_6_0_t183 = FSM_fft_64_stage_6_0_t182[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t184 = i_data_in_real[FSM_fft_64_stage_6_0_t183 * 32 +: 32];
    FSM_fft_64_stage_6_0_t185 = 32'b00000000000000000000000000101001;
    FSM_fft_64_stage_6_0_t186 = FSM_fft_64_stage_6_0_t185[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t187 = i_data_in_real[FSM_fft_64_stage_6_0_t186 * 32 +: 32];
    FSM_fft_64_stage_6_0_t188 = FSM_fft_64_stage_6_0_t184 + FSM_fft_64_stage_6_0_t187;
    FSM_fft_64_stage_6_0_t189 = FSM_fft_64_stage_6_0_t188[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t190 = FSM_fft_64_stage_6_0_t179;
    FSM_fft_64_stage_6_0_t190[FSM_fft_64_stage_6_0_t181 * 32 +: 32] = FSM_fft_64_stage_6_0_t189;
    FSM_fft_64_stage_6_0_t191 = 32'b00000000000000000000000000101001;
    FSM_fft_64_stage_6_0_t192 = FSM_fft_64_stage_6_0_t191[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t193 = 32'b00000000000000000000000000001001;
    FSM_fft_64_stage_6_0_t194 = FSM_fft_64_stage_6_0_t193[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t195 = i_data_in_real[FSM_fft_64_stage_6_0_t194 * 32 +: 32];
    FSM_fft_64_stage_6_0_t196 = 32'b00000000000000000000000000101001;
    FSM_fft_64_stage_6_0_t197 = FSM_fft_64_stage_6_0_t196[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t198 = i_data_in_real[FSM_fft_64_stage_6_0_t197 * 32 +: 32];
    FSM_fft_64_stage_6_0_t199 = FSM_fft_64_stage_6_0_t190;
    FSM_fft_64_stage_6_0_t199[FSM_fft_64_stage_6_0_t192 * 32 +: 32] = FSM_fft_64_stage_6_0_t195 - FSM_fft_64_stage_6_0_t198;
    FSM_fft_64_stage_6_0_t200 = 32'b00000000000000000000000000001010;
    FSM_fft_64_stage_6_0_t201 = FSM_fft_64_stage_6_0_t200[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t202 = 32'b00000000000000000000000000001010;
    FSM_fft_64_stage_6_0_t203 = FSM_fft_64_stage_6_0_t202[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t204 = i_data_in_real[FSM_fft_64_stage_6_0_t203 * 32 +: 32];
    FSM_fft_64_stage_6_0_t205 = 32'b00000000000000000000000000101010;
    FSM_fft_64_stage_6_0_t206 = FSM_fft_64_stage_6_0_t205[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t207 = i_data_in_real[FSM_fft_64_stage_6_0_t206 * 32 +: 32];
    FSM_fft_64_stage_6_0_t208 = FSM_fft_64_stage_6_0_t204 + FSM_fft_64_stage_6_0_t207;
    FSM_fft_64_stage_6_0_t209 = FSM_fft_64_stage_6_0_t208[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t210 = FSM_fft_64_stage_6_0_t199;
    FSM_fft_64_stage_6_0_t210[FSM_fft_64_stage_6_0_t201 * 32 +: 32] = FSM_fft_64_stage_6_0_t209;
    FSM_fft_64_stage_6_0_t211 = 32'b00000000000000000000000000101010;
    FSM_fft_64_stage_6_0_t212 = FSM_fft_64_stage_6_0_t211[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t213 = 32'b00000000000000000000000000001010;
    FSM_fft_64_stage_6_0_t214 = FSM_fft_64_stage_6_0_t213[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t215 = i_data_in_real[FSM_fft_64_stage_6_0_t214 * 32 +: 32];
    FSM_fft_64_stage_6_0_t216 = 32'b00000000000000000000000000101010;
    FSM_fft_64_stage_6_0_t217 = FSM_fft_64_stage_6_0_t216[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t218 = i_data_in_real[FSM_fft_64_stage_6_0_t217 * 32 +: 32];
    FSM_fft_64_stage_6_0_t219 = FSM_fft_64_stage_6_0_t210;
    FSM_fft_64_stage_6_0_t219[FSM_fft_64_stage_6_0_t212 * 32 +: 32] = FSM_fft_64_stage_6_0_t215 - FSM_fft_64_stage_6_0_t218;
    FSM_fft_64_stage_6_0_t220 = 32'b00000000000000000000000000001011;
    FSM_fft_64_stage_6_0_t221 = FSM_fft_64_stage_6_0_t220[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t222 = 32'b00000000000000000000000000001011;
    FSM_fft_64_stage_6_0_t223 = FSM_fft_64_stage_6_0_t222[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t224 = i_data_in_real[FSM_fft_64_stage_6_0_t223 * 32 +: 32];
    FSM_fft_64_stage_6_0_t225 = 32'b00000000000000000000000000101011;
    FSM_fft_64_stage_6_0_t226 = FSM_fft_64_stage_6_0_t225[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t227 = i_data_in_real[FSM_fft_64_stage_6_0_t226 * 32 +: 32];
    FSM_fft_64_stage_6_0_t228 = FSM_fft_64_stage_6_0_t224 + FSM_fft_64_stage_6_0_t227;
    FSM_fft_64_stage_6_0_t229 = FSM_fft_64_stage_6_0_t228[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t230 = FSM_fft_64_stage_6_0_t219;
    FSM_fft_64_stage_6_0_t230[FSM_fft_64_stage_6_0_t221 * 32 +: 32] = FSM_fft_64_stage_6_0_t229;
    FSM_fft_64_stage_6_0_t231 = 32'b00000000000000000000000000101011;
    FSM_fft_64_stage_6_0_t232 = FSM_fft_64_stage_6_0_t231[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t233 = 32'b00000000000000000000000000001011;
    FSM_fft_64_stage_6_0_t234 = FSM_fft_64_stage_6_0_t233[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t235 = i_data_in_real[FSM_fft_64_stage_6_0_t234 * 32 +: 32];
    FSM_fft_64_stage_6_0_t236 = 32'b00000000000000000000000000101011;
    FSM_fft_64_stage_6_0_t237 = FSM_fft_64_stage_6_0_t236[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t238 = i_data_in_real[FSM_fft_64_stage_6_0_t237 * 32 +: 32];
    FSM_fft_64_stage_6_0_t239 = FSM_fft_64_stage_6_0_t230;
    FSM_fft_64_stage_6_0_t239[FSM_fft_64_stage_6_0_t232 * 32 +: 32] = FSM_fft_64_stage_6_0_t235 - FSM_fft_64_stage_6_0_t238;
    FSM_fft_64_stage_6_0_t240 = 32'b00000000000000000000000000001100;
    FSM_fft_64_stage_6_0_t241 = FSM_fft_64_stage_6_0_t240[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t242 = 32'b00000000000000000000000000001100;
    FSM_fft_64_stage_6_0_t243 = FSM_fft_64_stage_6_0_t242[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t244 = i_data_in_real[FSM_fft_64_stage_6_0_t243 * 32 +: 32];
    FSM_fft_64_stage_6_0_t245 = 32'b00000000000000000000000000101100;
    FSM_fft_64_stage_6_0_t246 = FSM_fft_64_stage_6_0_t245[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t247 = i_data_in_real[FSM_fft_64_stage_6_0_t246 * 32 +: 32];
    FSM_fft_64_stage_6_0_t248 = FSM_fft_64_stage_6_0_t244 + FSM_fft_64_stage_6_0_t247;
    FSM_fft_64_stage_6_0_t249 = FSM_fft_64_stage_6_0_t248[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t250 = FSM_fft_64_stage_6_0_t239;
    FSM_fft_64_stage_6_0_t250[FSM_fft_64_stage_6_0_t241 * 32 +: 32] = FSM_fft_64_stage_6_0_t249;
    FSM_fft_64_stage_6_0_t251 = 32'b00000000000000000000000000101100;
    FSM_fft_64_stage_6_0_t252 = FSM_fft_64_stage_6_0_t251[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t253 = 32'b00000000000000000000000000001100;
    FSM_fft_64_stage_6_0_t254 = FSM_fft_64_stage_6_0_t253[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t255 = i_data_in_real[FSM_fft_64_stage_6_0_t254 * 32 +: 32];
    FSM_fft_64_stage_6_0_t256 = 32'b00000000000000000000000000101100;
    FSM_fft_64_stage_6_0_t257 = FSM_fft_64_stage_6_0_t256[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t258 = i_data_in_real[FSM_fft_64_stage_6_0_t257 * 32 +: 32];
    FSM_fft_64_stage_6_0_t259 = FSM_fft_64_stage_6_0_t250;
    FSM_fft_64_stage_6_0_t259[FSM_fft_64_stage_6_0_t252 * 32 +: 32] = FSM_fft_64_stage_6_0_t255 - FSM_fft_64_stage_6_0_t258;
    FSM_fft_64_stage_6_0_t260 = 32'b00000000000000000000000000001101;
    FSM_fft_64_stage_6_0_t261 = FSM_fft_64_stage_6_0_t260[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t262 = 32'b00000000000000000000000000001101;
    FSM_fft_64_stage_6_0_t263 = FSM_fft_64_stage_6_0_t262[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t264 = i_data_in_real[FSM_fft_64_stage_6_0_t263 * 32 +: 32];
    FSM_fft_64_stage_6_0_t265 = 32'b00000000000000000000000000101101;
    FSM_fft_64_stage_6_0_t266 = FSM_fft_64_stage_6_0_t265[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t267 = i_data_in_real[FSM_fft_64_stage_6_0_t266 * 32 +: 32];
    FSM_fft_64_stage_6_0_t268 = FSM_fft_64_stage_6_0_t264 + FSM_fft_64_stage_6_0_t267;
    FSM_fft_64_stage_6_0_t269 = FSM_fft_64_stage_6_0_t268[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t270 = FSM_fft_64_stage_6_0_t259;
    FSM_fft_64_stage_6_0_t270[FSM_fft_64_stage_6_0_t261 * 32 +: 32] = FSM_fft_64_stage_6_0_t269;
    FSM_fft_64_stage_6_0_t271 = 32'b00000000000000000000000000101101;
    FSM_fft_64_stage_6_0_t272 = FSM_fft_64_stage_6_0_t271[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t273 = 32'b00000000000000000000000000001101;
    FSM_fft_64_stage_6_0_t274 = FSM_fft_64_stage_6_0_t273[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t275 = i_data_in_real[FSM_fft_64_stage_6_0_t274 * 32 +: 32];
    FSM_fft_64_stage_6_0_t276 = 32'b00000000000000000000000000101101;
    FSM_fft_64_stage_6_0_t277 = FSM_fft_64_stage_6_0_t276[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t278 = i_data_in_real[FSM_fft_64_stage_6_0_t277 * 32 +: 32];
    FSM_fft_64_stage_6_0_t279 = FSM_fft_64_stage_6_0_t270;
    FSM_fft_64_stage_6_0_t279[FSM_fft_64_stage_6_0_t272 * 32 +: 32] = FSM_fft_64_stage_6_0_t275 - FSM_fft_64_stage_6_0_t278;
    FSM_fft_64_stage_6_0_t280 = 32'b00000000000000000000000000001110;
    FSM_fft_64_stage_6_0_t281 = FSM_fft_64_stage_6_0_t280[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t282 = 32'b00000000000000000000000000001110;
    FSM_fft_64_stage_6_0_t283 = FSM_fft_64_stage_6_0_t282[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t284 = i_data_in_real[FSM_fft_64_stage_6_0_t283 * 32 +: 32];
    FSM_fft_64_stage_6_0_t285 = 32'b00000000000000000000000000101110;
    FSM_fft_64_stage_6_0_t286 = FSM_fft_64_stage_6_0_t285[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t287 = i_data_in_real[FSM_fft_64_stage_6_0_t286 * 32 +: 32];
    FSM_fft_64_stage_6_0_t288 = FSM_fft_64_stage_6_0_t284 + FSM_fft_64_stage_6_0_t287;
    FSM_fft_64_stage_6_0_t289 = FSM_fft_64_stage_6_0_t288[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t290 = FSM_fft_64_stage_6_0_t279;
    FSM_fft_64_stage_6_0_t290[FSM_fft_64_stage_6_0_t281 * 32 +: 32] = FSM_fft_64_stage_6_0_t289;
    FSM_fft_64_stage_6_0_t291 = 32'b00000000000000000000000000101110;
    FSM_fft_64_stage_6_0_t292 = FSM_fft_64_stage_6_0_t291[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t293 = 32'b00000000000000000000000000001110;
    FSM_fft_64_stage_6_0_t294 = FSM_fft_64_stage_6_0_t293[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t295 = i_data_in_real[FSM_fft_64_stage_6_0_t294 * 32 +: 32];
    FSM_fft_64_stage_6_0_t296 = 32'b00000000000000000000000000101110;
    FSM_fft_64_stage_6_0_t297 = FSM_fft_64_stage_6_0_t296[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t298 = i_data_in_real[FSM_fft_64_stage_6_0_t297 * 32 +: 32];
    FSM_fft_64_stage_6_0_t299 = FSM_fft_64_stage_6_0_t290;
    FSM_fft_64_stage_6_0_t299[FSM_fft_64_stage_6_0_t292 * 32 +: 32] = FSM_fft_64_stage_6_0_t295 - FSM_fft_64_stage_6_0_t298;
    FSM_fft_64_stage_6_0_t300 = 32'b00000000000000000000000000001111;
    FSM_fft_64_stage_6_0_t301 = FSM_fft_64_stage_6_0_t300[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t302 = 32'b00000000000000000000000000001111;
    FSM_fft_64_stage_6_0_t303 = FSM_fft_64_stage_6_0_t302[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t304 = i_data_in_real[FSM_fft_64_stage_6_0_t303 * 32 +: 32];
    FSM_fft_64_stage_6_0_t305 = 32'b00000000000000000000000000101111;
    FSM_fft_64_stage_6_0_t306 = FSM_fft_64_stage_6_0_t305[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t307 = i_data_in_real[FSM_fft_64_stage_6_0_t306 * 32 +: 32];
    FSM_fft_64_stage_6_0_t308 = FSM_fft_64_stage_6_0_t304 + FSM_fft_64_stage_6_0_t307;
    FSM_fft_64_stage_6_0_t309 = FSM_fft_64_stage_6_0_t308[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t310 = FSM_fft_64_stage_6_0_t299;
    FSM_fft_64_stage_6_0_t310[FSM_fft_64_stage_6_0_t301 * 32 +: 32] = FSM_fft_64_stage_6_0_t309;
    FSM_fft_64_stage_6_0_t311 = 32'b00000000000000000000000000101111;
    FSM_fft_64_stage_6_0_t312 = FSM_fft_64_stage_6_0_t311[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t313 = 32'b00000000000000000000000000001111;
    FSM_fft_64_stage_6_0_t314 = FSM_fft_64_stage_6_0_t313[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t315 = i_data_in_real[FSM_fft_64_stage_6_0_t314 * 32 +: 32];
    FSM_fft_64_stage_6_0_t316 = 32'b00000000000000000000000000101111;
    FSM_fft_64_stage_6_0_t317 = FSM_fft_64_stage_6_0_t316[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t318 = i_data_in_real[FSM_fft_64_stage_6_0_t317 * 32 +: 32];
    FSM_fft_64_stage_6_0_t319 = FSM_fft_64_stage_6_0_t310;
    FSM_fft_64_stage_6_0_t319[FSM_fft_64_stage_6_0_t312 * 32 +: 32] = FSM_fft_64_stage_6_0_t315 - FSM_fft_64_stage_6_0_t318;
    FSM_fft_64_stage_6_0_t320 = 32'b00000000000000000000000000010000;
    FSM_fft_64_stage_6_0_t321 = FSM_fft_64_stage_6_0_t320[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t322 = 32'b00000000000000000000000000010000;
    FSM_fft_64_stage_6_0_t323 = FSM_fft_64_stage_6_0_t322[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t324 = i_data_in_real[FSM_fft_64_stage_6_0_t323 * 32 +: 32];
    FSM_fft_64_stage_6_0_t325 = 32'b00000000000000000000000000110000;
    FSM_fft_64_stage_6_0_t326 = FSM_fft_64_stage_6_0_t325[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t327 = i_data_in_real[FSM_fft_64_stage_6_0_t326 * 32 +: 32];
    FSM_fft_64_stage_6_0_t328 = FSM_fft_64_stage_6_0_t324 + FSM_fft_64_stage_6_0_t327;
    FSM_fft_64_stage_6_0_t329 = FSM_fft_64_stage_6_0_t328[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t330 = FSM_fft_64_stage_6_0_t319;
    FSM_fft_64_stage_6_0_t330[FSM_fft_64_stage_6_0_t321 * 32 +: 32] = FSM_fft_64_stage_6_0_t329;
    FSM_fft_64_stage_6_0_t331 = 32'b00000000000000000000000000110000;
    FSM_fft_64_stage_6_0_t332 = FSM_fft_64_stage_6_0_t331[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t333 = 32'b00000000000000000000000000010000;
    FSM_fft_64_stage_6_0_t334 = FSM_fft_64_stage_6_0_t333[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t335 = i_data_in_real[FSM_fft_64_stage_6_0_t334 * 32 +: 32];
    FSM_fft_64_stage_6_0_t336 = 32'b00000000000000000000000000110000;
    FSM_fft_64_stage_6_0_t337 = FSM_fft_64_stage_6_0_t336[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t338 = i_data_in_real[FSM_fft_64_stage_6_0_t337 * 32 +: 32];
    FSM_fft_64_stage_6_0_t339 = FSM_fft_64_stage_6_0_t330;
    FSM_fft_64_stage_6_0_t339[FSM_fft_64_stage_6_0_t332 * 32 +: 32] = FSM_fft_64_stage_6_0_t335 - FSM_fft_64_stage_6_0_t338;
    FSM_fft_64_stage_6_0_t340 = 32'b00000000000000000000000000010001;
    FSM_fft_64_stage_6_0_t341 = FSM_fft_64_stage_6_0_t340[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t342 = 32'b00000000000000000000000000010001;
    FSM_fft_64_stage_6_0_t343 = FSM_fft_64_stage_6_0_t342[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t344 = i_data_in_real[FSM_fft_64_stage_6_0_t343 * 32 +: 32];
    FSM_fft_64_stage_6_0_t345 = 32'b00000000000000000000000000110001;
    FSM_fft_64_stage_6_0_t346 = FSM_fft_64_stage_6_0_t345[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t347 = i_data_in_real[FSM_fft_64_stage_6_0_t346 * 32 +: 32];
    FSM_fft_64_stage_6_0_t348 = FSM_fft_64_stage_6_0_t344 + FSM_fft_64_stage_6_0_t347;
    FSM_fft_64_stage_6_0_t349 = FSM_fft_64_stage_6_0_t348[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t350 = FSM_fft_64_stage_6_0_t339;
    FSM_fft_64_stage_6_0_t350[FSM_fft_64_stage_6_0_t341 * 32 +: 32] = FSM_fft_64_stage_6_0_t349;
    FSM_fft_64_stage_6_0_t351 = 32'b00000000000000000000000000110001;
    FSM_fft_64_stage_6_0_t352 = FSM_fft_64_stage_6_0_t351[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t353 = 32'b00000000000000000000000000010001;
    FSM_fft_64_stage_6_0_t354 = FSM_fft_64_stage_6_0_t353[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t355 = i_data_in_real[FSM_fft_64_stage_6_0_t354 * 32 +: 32];
    FSM_fft_64_stage_6_0_t356 = 32'b00000000000000000000000000110001;
    FSM_fft_64_stage_6_0_t357 = FSM_fft_64_stage_6_0_t356[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t358 = i_data_in_real[FSM_fft_64_stage_6_0_t357 * 32 +: 32];
    FSM_fft_64_stage_6_0_t359 = FSM_fft_64_stage_6_0_t350;
    FSM_fft_64_stage_6_0_t359[FSM_fft_64_stage_6_0_t352 * 32 +: 32] = FSM_fft_64_stage_6_0_t355 - FSM_fft_64_stage_6_0_t358;
    FSM_fft_64_stage_6_0_t360 = 32'b00000000000000000000000000010010;
    FSM_fft_64_stage_6_0_t361 = FSM_fft_64_stage_6_0_t360[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t362 = 32'b00000000000000000000000000010010;
    FSM_fft_64_stage_6_0_t363 = FSM_fft_64_stage_6_0_t362[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t364 = i_data_in_real[FSM_fft_64_stage_6_0_t363 * 32 +: 32];
    FSM_fft_64_stage_6_0_t365 = 32'b00000000000000000000000000110010;
    FSM_fft_64_stage_6_0_t366 = FSM_fft_64_stage_6_0_t365[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t367 = i_data_in_real[FSM_fft_64_stage_6_0_t366 * 32 +: 32];
    FSM_fft_64_stage_6_0_t368 = FSM_fft_64_stage_6_0_t364 + FSM_fft_64_stage_6_0_t367;
    FSM_fft_64_stage_6_0_t369 = FSM_fft_64_stage_6_0_t368[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t370 = FSM_fft_64_stage_6_0_t359;
    FSM_fft_64_stage_6_0_t370[FSM_fft_64_stage_6_0_t361 * 32 +: 32] = FSM_fft_64_stage_6_0_t369;
    FSM_fft_64_stage_6_0_t371 = 32'b00000000000000000000000000110010;
    FSM_fft_64_stage_6_0_t372 = FSM_fft_64_stage_6_0_t371[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t373 = 32'b00000000000000000000000000010010;
    FSM_fft_64_stage_6_0_t374 = FSM_fft_64_stage_6_0_t373[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t375 = i_data_in_real[FSM_fft_64_stage_6_0_t374 * 32 +: 32];
    FSM_fft_64_stage_6_0_t376 = 32'b00000000000000000000000000110010;
    FSM_fft_64_stage_6_0_t377 = FSM_fft_64_stage_6_0_t376[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t378 = i_data_in_real[FSM_fft_64_stage_6_0_t377 * 32 +: 32];
    FSM_fft_64_stage_6_0_t379 = FSM_fft_64_stage_6_0_t370;
    FSM_fft_64_stage_6_0_t379[FSM_fft_64_stage_6_0_t372 * 32 +: 32] = FSM_fft_64_stage_6_0_t375 - FSM_fft_64_stage_6_0_t378;
    FSM_fft_64_stage_6_0_t380 = 32'b00000000000000000000000000010011;
    FSM_fft_64_stage_6_0_t381 = FSM_fft_64_stage_6_0_t380[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t382 = 32'b00000000000000000000000000010011;
    FSM_fft_64_stage_6_0_t383 = FSM_fft_64_stage_6_0_t382[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t384 = i_data_in_real[FSM_fft_64_stage_6_0_t383 * 32 +: 32];
    FSM_fft_64_stage_6_0_t385 = 32'b00000000000000000000000000110011;
    FSM_fft_64_stage_6_0_t386 = FSM_fft_64_stage_6_0_t385[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t387 = i_data_in_real[FSM_fft_64_stage_6_0_t386 * 32 +: 32];
    FSM_fft_64_stage_6_0_t388 = FSM_fft_64_stage_6_0_t384 + FSM_fft_64_stage_6_0_t387;
    FSM_fft_64_stage_6_0_t389 = FSM_fft_64_stage_6_0_t388[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t390 = FSM_fft_64_stage_6_0_t379;
    FSM_fft_64_stage_6_0_t390[FSM_fft_64_stage_6_0_t381 * 32 +: 32] = FSM_fft_64_stage_6_0_t389;
    FSM_fft_64_stage_6_0_t391 = 32'b00000000000000000000000000110011;
    FSM_fft_64_stage_6_0_t392 = FSM_fft_64_stage_6_0_t391[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t393 = 32'b00000000000000000000000000010011;
    FSM_fft_64_stage_6_0_t394 = FSM_fft_64_stage_6_0_t393[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t395 = i_data_in_real[FSM_fft_64_stage_6_0_t394 * 32 +: 32];
    FSM_fft_64_stage_6_0_t396 = 32'b00000000000000000000000000110011;
    FSM_fft_64_stage_6_0_t397 = FSM_fft_64_stage_6_0_t396[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t398 = i_data_in_real[FSM_fft_64_stage_6_0_t397 * 32 +: 32];
    FSM_fft_64_stage_6_0_t399 = FSM_fft_64_stage_6_0_t390;
    FSM_fft_64_stage_6_0_t399[FSM_fft_64_stage_6_0_t392 * 32 +: 32] = FSM_fft_64_stage_6_0_t395 - FSM_fft_64_stage_6_0_t398;
    FSM_fft_64_stage_6_0_t400 = 32'b00000000000000000000000000010100;
    FSM_fft_64_stage_6_0_t401 = FSM_fft_64_stage_6_0_t400[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t402 = 32'b00000000000000000000000000010100;
    FSM_fft_64_stage_6_0_t403 = FSM_fft_64_stage_6_0_t402[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t404 = i_data_in_real[FSM_fft_64_stage_6_0_t403 * 32 +: 32];
    FSM_fft_64_stage_6_0_t405 = 32'b00000000000000000000000000110100;
    FSM_fft_64_stage_6_0_t406 = FSM_fft_64_stage_6_0_t405[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t407 = i_data_in_real[FSM_fft_64_stage_6_0_t406 * 32 +: 32];
    FSM_fft_64_stage_6_0_t408 = FSM_fft_64_stage_6_0_t404 + FSM_fft_64_stage_6_0_t407;
    FSM_fft_64_stage_6_0_t409 = FSM_fft_64_stage_6_0_t408[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t410 = FSM_fft_64_stage_6_0_t399;
    FSM_fft_64_stage_6_0_t410[FSM_fft_64_stage_6_0_t401 * 32 +: 32] = FSM_fft_64_stage_6_0_t409;
    FSM_fft_64_stage_6_0_t411 = 32'b00000000000000000000000000110100;
    FSM_fft_64_stage_6_0_t412 = FSM_fft_64_stage_6_0_t411[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t413 = 32'b00000000000000000000000000010100;
    FSM_fft_64_stage_6_0_t414 = FSM_fft_64_stage_6_0_t413[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t415 = i_data_in_real[FSM_fft_64_stage_6_0_t414 * 32 +: 32];
    FSM_fft_64_stage_6_0_t416 = 32'b00000000000000000000000000110100;
    FSM_fft_64_stage_6_0_t417 = FSM_fft_64_stage_6_0_t416[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t418 = i_data_in_real[FSM_fft_64_stage_6_0_t417 * 32 +: 32];
    FSM_fft_64_stage_6_0_t419 = FSM_fft_64_stage_6_0_t410;
    FSM_fft_64_stage_6_0_t419[FSM_fft_64_stage_6_0_t412 * 32 +: 32] = FSM_fft_64_stage_6_0_t415 - FSM_fft_64_stage_6_0_t418;
    FSM_fft_64_stage_6_0_t420 = 32'b00000000000000000000000000010101;
    FSM_fft_64_stage_6_0_t421 = FSM_fft_64_stage_6_0_t420[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t422 = 32'b00000000000000000000000000010101;
    FSM_fft_64_stage_6_0_t423 = FSM_fft_64_stage_6_0_t422[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t424 = i_data_in_real[FSM_fft_64_stage_6_0_t423 * 32 +: 32];
    FSM_fft_64_stage_6_0_t425 = 32'b00000000000000000000000000110101;
    FSM_fft_64_stage_6_0_t426 = FSM_fft_64_stage_6_0_t425[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t427 = i_data_in_real[FSM_fft_64_stage_6_0_t426 * 32 +: 32];
    FSM_fft_64_stage_6_0_t428 = FSM_fft_64_stage_6_0_t424 + FSM_fft_64_stage_6_0_t427;
    FSM_fft_64_stage_6_0_t429 = FSM_fft_64_stage_6_0_t428[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t430 = FSM_fft_64_stage_6_0_t419;
    FSM_fft_64_stage_6_0_t430[FSM_fft_64_stage_6_0_t421 * 32 +: 32] = FSM_fft_64_stage_6_0_t429;
    FSM_fft_64_stage_6_0_t431 = 32'b00000000000000000000000000110101;
    FSM_fft_64_stage_6_0_t432 = FSM_fft_64_stage_6_0_t431[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t433 = 32'b00000000000000000000000000010101;
    FSM_fft_64_stage_6_0_t434 = FSM_fft_64_stage_6_0_t433[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t435 = i_data_in_real[FSM_fft_64_stage_6_0_t434 * 32 +: 32];
    FSM_fft_64_stage_6_0_t436 = 32'b00000000000000000000000000110101;
    FSM_fft_64_stage_6_0_t437 = FSM_fft_64_stage_6_0_t436[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t438 = i_data_in_real[FSM_fft_64_stage_6_0_t437 * 32 +: 32];
    FSM_fft_64_stage_6_0_t439 = FSM_fft_64_stage_6_0_t430;
    FSM_fft_64_stage_6_0_t439[FSM_fft_64_stage_6_0_t432 * 32 +: 32] = FSM_fft_64_stage_6_0_t435 - FSM_fft_64_stage_6_0_t438;
    FSM_fft_64_stage_6_0_t440 = 32'b00000000000000000000000000010110;
    FSM_fft_64_stage_6_0_t441 = FSM_fft_64_stage_6_0_t440[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t442 = 32'b00000000000000000000000000010110;
    FSM_fft_64_stage_6_0_t443 = FSM_fft_64_stage_6_0_t442[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t444 = i_data_in_real[FSM_fft_64_stage_6_0_t443 * 32 +: 32];
    FSM_fft_64_stage_6_0_t445 = 32'b00000000000000000000000000110110;
    FSM_fft_64_stage_6_0_t446 = FSM_fft_64_stage_6_0_t445[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t447 = i_data_in_real[FSM_fft_64_stage_6_0_t446 * 32 +: 32];
    FSM_fft_64_stage_6_0_t448 = FSM_fft_64_stage_6_0_t444 + FSM_fft_64_stage_6_0_t447;
    FSM_fft_64_stage_6_0_t449 = FSM_fft_64_stage_6_0_t448[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t450 = FSM_fft_64_stage_6_0_t439;
    FSM_fft_64_stage_6_0_t450[FSM_fft_64_stage_6_0_t441 * 32 +: 32] = FSM_fft_64_stage_6_0_t449;
    FSM_fft_64_stage_6_0_t451 = 32'b00000000000000000000000000110110;
    FSM_fft_64_stage_6_0_t452 = FSM_fft_64_stage_6_0_t451[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t453 = 32'b00000000000000000000000000010110;
    FSM_fft_64_stage_6_0_t454 = FSM_fft_64_stage_6_0_t453[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t455 = i_data_in_real[FSM_fft_64_stage_6_0_t454 * 32 +: 32];
    FSM_fft_64_stage_6_0_t456 = 32'b00000000000000000000000000110110;
    FSM_fft_64_stage_6_0_t457 = FSM_fft_64_stage_6_0_t456[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t458 = i_data_in_real[FSM_fft_64_stage_6_0_t457 * 32 +: 32];
    FSM_fft_64_stage_6_0_t459 = FSM_fft_64_stage_6_0_t450;
    FSM_fft_64_stage_6_0_t459[FSM_fft_64_stage_6_0_t452 * 32 +: 32] = FSM_fft_64_stage_6_0_t455 - FSM_fft_64_stage_6_0_t458;
    FSM_fft_64_stage_6_0_t460 = 32'b00000000000000000000000000010111;
    FSM_fft_64_stage_6_0_t461 = FSM_fft_64_stage_6_0_t460[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t462 = 32'b00000000000000000000000000010111;
    FSM_fft_64_stage_6_0_t463 = FSM_fft_64_stage_6_0_t462[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t464 = i_data_in_real[FSM_fft_64_stage_6_0_t463 * 32 +: 32];
    FSM_fft_64_stage_6_0_t465 = 32'b00000000000000000000000000110111;
    FSM_fft_64_stage_6_0_t466 = FSM_fft_64_stage_6_0_t465[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t467 = i_data_in_real[FSM_fft_64_stage_6_0_t466 * 32 +: 32];
    FSM_fft_64_stage_6_0_t468 = FSM_fft_64_stage_6_0_t464 + FSM_fft_64_stage_6_0_t467;
    FSM_fft_64_stage_6_0_t469 = FSM_fft_64_stage_6_0_t468[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t470 = FSM_fft_64_stage_6_0_t459;
    FSM_fft_64_stage_6_0_t470[FSM_fft_64_stage_6_0_t461 * 32 +: 32] = FSM_fft_64_stage_6_0_t469;
    FSM_fft_64_stage_6_0_t471 = 32'b00000000000000000000000000110111;
    FSM_fft_64_stage_6_0_t472 = FSM_fft_64_stage_6_0_t471[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t473 = 32'b00000000000000000000000000010111;
    FSM_fft_64_stage_6_0_t474 = FSM_fft_64_stage_6_0_t473[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t475 = i_data_in_real[FSM_fft_64_stage_6_0_t474 * 32 +: 32];
    FSM_fft_64_stage_6_0_t476 = 32'b00000000000000000000000000110111;
    FSM_fft_64_stage_6_0_t477 = FSM_fft_64_stage_6_0_t476[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t478 = i_data_in_real[FSM_fft_64_stage_6_0_t477 * 32 +: 32];
    FSM_fft_64_stage_6_0_t479 = FSM_fft_64_stage_6_0_t470;
    FSM_fft_64_stage_6_0_t479[FSM_fft_64_stage_6_0_t472 * 32 +: 32] = FSM_fft_64_stage_6_0_t475 - FSM_fft_64_stage_6_0_t478;
    FSM_fft_64_stage_6_0_t480 = 32'b00000000000000000000000000011000;
    FSM_fft_64_stage_6_0_t481 = FSM_fft_64_stage_6_0_t480[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t482 = 32'b00000000000000000000000000011000;
    FSM_fft_64_stage_6_0_t483 = FSM_fft_64_stage_6_0_t482[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t484 = i_data_in_real[FSM_fft_64_stage_6_0_t483 * 32 +: 32];
    FSM_fft_64_stage_6_0_t485 = 32'b00000000000000000000000000111000;
    FSM_fft_64_stage_6_0_t486 = FSM_fft_64_stage_6_0_t485[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t487 = i_data_in_real[FSM_fft_64_stage_6_0_t486 * 32 +: 32];
    FSM_fft_64_stage_6_0_t488 = FSM_fft_64_stage_6_0_t484 + FSM_fft_64_stage_6_0_t487;
    FSM_fft_64_stage_6_0_t489 = FSM_fft_64_stage_6_0_t488[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t490 = FSM_fft_64_stage_6_0_t479;
    FSM_fft_64_stage_6_0_t490[FSM_fft_64_stage_6_0_t481 * 32 +: 32] = FSM_fft_64_stage_6_0_t489;
    FSM_fft_64_stage_6_0_t491 = 32'b00000000000000000000000000111000;
    FSM_fft_64_stage_6_0_t492 = FSM_fft_64_stage_6_0_t491[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t493 = 32'b00000000000000000000000000011000;
    FSM_fft_64_stage_6_0_t494 = FSM_fft_64_stage_6_0_t493[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t495 = i_data_in_real[FSM_fft_64_stage_6_0_t494 * 32 +: 32];
    FSM_fft_64_stage_6_0_t496 = 32'b00000000000000000000000000111000;
    FSM_fft_64_stage_6_0_t497 = FSM_fft_64_stage_6_0_t496[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t498 = i_data_in_real[FSM_fft_64_stage_6_0_t497 * 32 +: 32];
    FSM_fft_64_stage_6_0_t499 = FSM_fft_64_stage_6_0_t490;
    FSM_fft_64_stage_6_0_t499[FSM_fft_64_stage_6_0_t492 * 32 +: 32] = FSM_fft_64_stage_6_0_t495 - FSM_fft_64_stage_6_0_t498;
    FSM_fft_64_stage_6_0_t500 = 32'b00000000000000000000000000011001;
    FSM_fft_64_stage_6_0_t501 = FSM_fft_64_stage_6_0_t500[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t502 = 32'b00000000000000000000000000011001;
    FSM_fft_64_stage_6_0_t503 = FSM_fft_64_stage_6_0_t502[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t504 = i_data_in_real[FSM_fft_64_stage_6_0_t503 * 32 +: 32];
    FSM_fft_64_stage_6_0_t505 = 32'b00000000000000000000000000111001;
    FSM_fft_64_stage_6_0_t506 = FSM_fft_64_stage_6_0_t505[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t507 = i_data_in_real[FSM_fft_64_stage_6_0_t506 * 32 +: 32];
    FSM_fft_64_stage_6_0_t508 = FSM_fft_64_stage_6_0_t504 + FSM_fft_64_stage_6_0_t507;
    FSM_fft_64_stage_6_0_t509 = FSM_fft_64_stage_6_0_t508[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t510 = FSM_fft_64_stage_6_0_t499;
    FSM_fft_64_stage_6_0_t510[FSM_fft_64_stage_6_0_t501 * 32 +: 32] = FSM_fft_64_stage_6_0_t509;
    FSM_fft_64_stage_6_0_t511 = 32'b00000000000000000000000000111001;
    FSM_fft_64_stage_6_0_t512 = FSM_fft_64_stage_6_0_t511[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t513 = 32'b00000000000000000000000000011001;
    FSM_fft_64_stage_6_0_t514 = FSM_fft_64_stage_6_0_t513[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t515 = i_data_in_real[FSM_fft_64_stage_6_0_t514 * 32 +: 32];
    FSM_fft_64_stage_6_0_t516 = 32'b00000000000000000000000000111001;
    FSM_fft_64_stage_6_0_t517 = FSM_fft_64_stage_6_0_t516[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t518 = i_data_in_real[FSM_fft_64_stage_6_0_t517 * 32 +: 32];
    FSM_fft_64_stage_6_0_t519 = FSM_fft_64_stage_6_0_t510;
    FSM_fft_64_stage_6_0_t519[FSM_fft_64_stage_6_0_t512 * 32 +: 32] = FSM_fft_64_stage_6_0_t515 - FSM_fft_64_stage_6_0_t518;
    FSM_fft_64_stage_6_0_t520 = 32'b00000000000000000000000000011010;
    FSM_fft_64_stage_6_0_t521 = FSM_fft_64_stage_6_0_t520[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t522 = 32'b00000000000000000000000000011010;
    FSM_fft_64_stage_6_0_t523 = FSM_fft_64_stage_6_0_t522[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t524 = i_data_in_real[FSM_fft_64_stage_6_0_t523 * 32 +: 32];
    FSM_fft_64_stage_6_0_t525 = 32'b00000000000000000000000000111010;
    FSM_fft_64_stage_6_0_t526 = FSM_fft_64_stage_6_0_t525[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t527 = i_data_in_real[FSM_fft_64_stage_6_0_t526 * 32 +: 32];
    FSM_fft_64_stage_6_0_t528 = FSM_fft_64_stage_6_0_t524 + FSM_fft_64_stage_6_0_t527;
    FSM_fft_64_stage_6_0_t529 = FSM_fft_64_stage_6_0_t528[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t530 = FSM_fft_64_stage_6_0_t519;
    FSM_fft_64_stage_6_0_t530[FSM_fft_64_stage_6_0_t521 * 32 +: 32] = FSM_fft_64_stage_6_0_t529;
    FSM_fft_64_stage_6_0_t531 = 32'b00000000000000000000000000111010;
    FSM_fft_64_stage_6_0_t532 = FSM_fft_64_stage_6_0_t531[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t533 = 32'b00000000000000000000000000011010;
    FSM_fft_64_stage_6_0_t534 = FSM_fft_64_stage_6_0_t533[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t535 = i_data_in_real[FSM_fft_64_stage_6_0_t534 * 32 +: 32];
    FSM_fft_64_stage_6_0_t536 = 32'b00000000000000000000000000111010;
    FSM_fft_64_stage_6_0_t537 = FSM_fft_64_stage_6_0_t536[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t538 = i_data_in_real[FSM_fft_64_stage_6_0_t537 * 32 +: 32];
    FSM_fft_64_stage_6_0_t539 = FSM_fft_64_stage_6_0_t530;
    FSM_fft_64_stage_6_0_t539[FSM_fft_64_stage_6_0_t532 * 32 +: 32] = FSM_fft_64_stage_6_0_t535 - FSM_fft_64_stage_6_0_t538;
    FSM_fft_64_stage_6_0_t540 = 32'b00000000000000000000000000011011;
    FSM_fft_64_stage_6_0_t541 = FSM_fft_64_stage_6_0_t540[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t542 = 32'b00000000000000000000000000011011;
    FSM_fft_64_stage_6_0_t543 = FSM_fft_64_stage_6_0_t542[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t544 = i_data_in_real[FSM_fft_64_stage_6_0_t543 * 32 +: 32];
    FSM_fft_64_stage_6_0_t545 = 32'b00000000000000000000000000111011;
    FSM_fft_64_stage_6_0_t546 = FSM_fft_64_stage_6_0_t545[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t547 = i_data_in_real[FSM_fft_64_stage_6_0_t546 * 32 +: 32];
    FSM_fft_64_stage_6_0_t548 = FSM_fft_64_stage_6_0_t544 + FSM_fft_64_stage_6_0_t547;
    FSM_fft_64_stage_6_0_t549 = FSM_fft_64_stage_6_0_t548[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t550 = FSM_fft_64_stage_6_0_t539;
    FSM_fft_64_stage_6_0_t550[FSM_fft_64_stage_6_0_t541 * 32 +: 32] = FSM_fft_64_stage_6_0_t549;
    FSM_fft_64_stage_6_0_t551 = 32'b00000000000000000000000000111011;
    FSM_fft_64_stage_6_0_t552 = FSM_fft_64_stage_6_0_t551[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t553 = 32'b00000000000000000000000000011011;
    FSM_fft_64_stage_6_0_t554 = FSM_fft_64_stage_6_0_t553[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t555 = i_data_in_real[FSM_fft_64_stage_6_0_t554 * 32 +: 32];
    FSM_fft_64_stage_6_0_t556 = 32'b00000000000000000000000000111011;
    FSM_fft_64_stage_6_0_t557 = FSM_fft_64_stage_6_0_t556[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t558 = i_data_in_real[FSM_fft_64_stage_6_0_t557 * 32 +: 32];
    FSM_fft_64_stage_6_0_t559 = FSM_fft_64_stage_6_0_t550;
    FSM_fft_64_stage_6_0_t559[FSM_fft_64_stage_6_0_t552 * 32 +: 32] = FSM_fft_64_stage_6_0_t555 - FSM_fft_64_stage_6_0_t558;
    FSM_fft_64_stage_6_0_t560 = 32'b00000000000000000000000000011100;
    FSM_fft_64_stage_6_0_t561 = FSM_fft_64_stage_6_0_t560[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t562 = 32'b00000000000000000000000000011100;
    FSM_fft_64_stage_6_0_t563 = FSM_fft_64_stage_6_0_t562[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t564 = i_data_in_real[FSM_fft_64_stage_6_0_t563 * 32 +: 32];
    FSM_fft_64_stage_6_0_t565 = 32'b00000000000000000000000000111100;
    FSM_fft_64_stage_6_0_t566 = FSM_fft_64_stage_6_0_t565[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t567 = i_data_in_real[FSM_fft_64_stage_6_0_t566 * 32 +: 32];
    FSM_fft_64_stage_6_0_t568 = FSM_fft_64_stage_6_0_t564 + FSM_fft_64_stage_6_0_t567;
    FSM_fft_64_stage_6_0_t569 = FSM_fft_64_stage_6_0_t568[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t570 = FSM_fft_64_stage_6_0_t559;
    FSM_fft_64_stage_6_0_t570[FSM_fft_64_stage_6_0_t561 * 32 +: 32] = FSM_fft_64_stage_6_0_t569;
    FSM_fft_64_stage_6_0_t571 = 32'b00000000000000000000000000111100;
    FSM_fft_64_stage_6_0_t572 = FSM_fft_64_stage_6_0_t571[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t573 = 32'b00000000000000000000000000011100;
    FSM_fft_64_stage_6_0_t574 = FSM_fft_64_stage_6_0_t573[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t575 = i_data_in_real[FSM_fft_64_stage_6_0_t574 * 32 +: 32];
    FSM_fft_64_stage_6_0_t576 = 32'b00000000000000000000000000111100;
    FSM_fft_64_stage_6_0_t577 = FSM_fft_64_stage_6_0_t576[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t578 = i_data_in_real[FSM_fft_64_stage_6_0_t577 * 32 +: 32];
    FSM_fft_64_stage_6_0_t579 = FSM_fft_64_stage_6_0_t570;
    FSM_fft_64_stage_6_0_t579[FSM_fft_64_stage_6_0_t572 * 32 +: 32] = FSM_fft_64_stage_6_0_t575 - FSM_fft_64_stage_6_0_t578;
    FSM_fft_64_stage_6_0_t580 = 32'b00000000000000000000000000011101;
    FSM_fft_64_stage_6_0_t581 = FSM_fft_64_stage_6_0_t580[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t582 = 32'b00000000000000000000000000011101;
    FSM_fft_64_stage_6_0_t583 = FSM_fft_64_stage_6_0_t582[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t584 = i_data_in_real[FSM_fft_64_stage_6_0_t583 * 32 +: 32];
    FSM_fft_64_stage_6_0_t585 = 32'b00000000000000000000000000111101;
    FSM_fft_64_stage_6_0_t586 = FSM_fft_64_stage_6_0_t585[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t587 = i_data_in_real[FSM_fft_64_stage_6_0_t586 * 32 +: 32];
    FSM_fft_64_stage_6_0_t588 = FSM_fft_64_stage_6_0_t584 + FSM_fft_64_stage_6_0_t587;
    FSM_fft_64_stage_6_0_t589 = FSM_fft_64_stage_6_0_t588[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t590 = FSM_fft_64_stage_6_0_t579;
    FSM_fft_64_stage_6_0_t590[FSM_fft_64_stage_6_0_t581 * 32 +: 32] = FSM_fft_64_stage_6_0_t589;
    FSM_fft_64_stage_6_0_t591 = 32'b00000000000000000000000000111101;
    FSM_fft_64_stage_6_0_t592 = FSM_fft_64_stage_6_0_t591[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t593 = 32'b00000000000000000000000000011101;
    FSM_fft_64_stage_6_0_t594 = FSM_fft_64_stage_6_0_t593[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t595 = i_data_in_real[FSM_fft_64_stage_6_0_t594 * 32 +: 32];
    FSM_fft_64_stage_6_0_t596 = 32'b00000000000000000000000000111101;
    FSM_fft_64_stage_6_0_t597 = FSM_fft_64_stage_6_0_t596[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t598 = i_data_in_real[FSM_fft_64_stage_6_0_t597 * 32 +: 32];
    FSM_fft_64_stage_6_0_t599 = FSM_fft_64_stage_6_0_t590;
    FSM_fft_64_stage_6_0_t599[FSM_fft_64_stage_6_0_t592 * 32 +: 32] = FSM_fft_64_stage_6_0_t595 - FSM_fft_64_stage_6_0_t598;
    FSM_fft_64_stage_6_0_t600 = 32'b00000000000000000000000000011110;
    FSM_fft_64_stage_6_0_t601 = FSM_fft_64_stage_6_0_t600[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t602 = 32'b00000000000000000000000000011110;
    FSM_fft_64_stage_6_0_t603 = FSM_fft_64_stage_6_0_t602[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t604 = i_data_in_real[FSM_fft_64_stage_6_0_t603 * 32 +: 32];
    FSM_fft_64_stage_6_0_t605 = 32'b00000000000000000000000000111110;
    FSM_fft_64_stage_6_0_t606 = FSM_fft_64_stage_6_0_t605[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t607 = i_data_in_real[FSM_fft_64_stage_6_0_t606 * 32 +: 32];
    FSM_fft_64_stage_6_0_t608 = FSM_fft_64_stage_6_0_t604 + FSM_fft_64_stage_6_0_t607;
    FSM_fft_64_stage_6_0_t609 = FSM_fft_64_stage_6_0_t608[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t610 = FSM_fft_64_stage_6_0_t599;
    FSM_fft_64_stage_6_0_t610[FSM_fft_64_stage_6_0_t601 * 32 +: 32] = FSM_fft_64_stage_6_0_t609;
    FSM_fft_64_stage_6_0_t611 = 32'b00000000000000000000000000111110;
    FSM_fft_64_stage_6_0_t612 = FSM_fft_64_stage_6_0_t611[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t613 = 32'b00000000000000000000000000011110;
    FSM_fft_64_stage_6_0_t614 = FSM_fft_64_stage_6_0_t613[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t615 = i_data_in_real[FSM_fft_64_stage_6_0_t614 * 32 +: 32];
    FSM_fft_64_stage_6_0_t616 = 32'b00000000000000000000000000111110;
    FSM_fft_64_stage_6_0_t617 = FSM_fft_64_stage_6_0_t616[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t618 = i_data_in_real[FSM_fft_64_stage_6_0_t617 * 32 +: 32];
    FSM_fft_64_stage_6_0_t619 = FSM_fft_64_stage_6_0_t610;
    FSM_fft_64_stage_6_0_t619[FSM_fft_64_stage_6_0_t612 * 32 +: 32] = FSM_fft_64_stage_6_0_t615 - FSM_fft_64_stage_6_0_t618;
    FSM_fft_64_stage_6_0_t620 = 32'b00000000000000000000000000011111;
    FSM_fft_64_stage_6_0_t621 = FSM_fft_64_stage_6_0_t620[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t622 = 32'b00000000000000000000000000011111;
    FSM_fft_64_stage_6_0_t623 = FSM_fft_64_stage_6_0_t622[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t624 = i_data_in_real[FSM_fft_64_stage_6_0_t623 * 32 +: 32];
    FSM_fft_64_stage_6_0_t625 = 32'b00000000000000000000000000111111;
    FSM_fft_64_stage_6_0_t626 = FSM_fft_64_stage_6_0_t625[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t627 = i_data_in_real[FSM_fft_64_stage_6_0_t626 * 32 +: 32];
    FSM_fft_64_stage_6_0_t628 = FSM_fft_64_stage_6_0_t624 + FSM_fft_64_stage_6_0_t627;
    FSM_fft_64_stage_6_0_t629 = FSM_fft_64_stage_6_0_t628[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t630 = FSM_fft_64_stage_6_0_t619;
    FSM_fft_64_stage_6_0_t630[FSM_fft_64_stage_6_0_t621 * 32 +: 32] = FSM_fft_64_stage_6_0_t629;
    FSM_fft_64_stage_6_0_t631 = 32'b00000000000000000000000000111111;
    FSM_fft_64_stage_6_0_t632 = FSM_fft_64_stage_6_0_t631[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t633 = 32'b00000000000000000000000000011111;
    FSM_fft_64_stage_6_0_t634 = FSM_fft_64_stage_6_0_t633[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t635 = i_data_in_real[FSM_fft_64_stage_6_0_t634 * 32 +: 32];
    FSM_fft_64_stage_6_0_t636 = 32'b00000000000000000000000000111111;
    FSM_fft_64_stage_6_0_t637 = FSM_fft_64_stage_6_0_t636[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t638 = i_data_in_real[FSM_fft_64_stage_6_0_t637 * 32 +: 32];
    FSM_fft_64_stage_6_0_t639 = FSM_fft_64_stage_6_0_t630;
    FSM_fft_64_stage_6_0_t639[FSM_fft_64_stage_6_0_t632 * 32 +: 32] = FSM_fft_64_stage_6_0_t635 - FSM_fft_64_stage_6_0_t638;
    FSM_fft_64_stage_6_0_t640 = 32'b0;
    FSM_fft_64_stage_6_0_t641 = FSM_fft_64_stage_6_0_t640[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t642 = 32'b0;
    FSM_fft_64_stage_6_0_t643 = FSM_fft_64_stage_6_0_t642[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t644 = i_data_in_imag[FSM_fft_64_stage_6_0_t643 * 32 +: 32];
    FSM_fft_64_stage_6_0_t645 = 32'b00000000000000000000000000100000;
    FSM_fft_64_stage_6_0_t646 = FSM_fft_64_stage_6_0_t645[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t647 = i_data_in_imag[FSM_fft_64_stage_6_0_t646 * 32 +: 32];
    FSM_fft_64_stage_6_0_t648 = FSM_fft_64_stage_6_0_t644 + FSM_fft_64_stage_6_0_t647;
    FSM_fft_64_stage_6_0_t649 = FSM_fft_64_stage_6_0_t648[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t650 = i_data_in_imag;
    FSM_fft_64_stage_6_0_t650[FSM_fft_64_stage_6_0_t641 * 32 +: 32] = FSM_fft_64_stage_6_0_t649;
    FSM_fft_64_stage_6_0_t651 = 32'b00000000000000000000000000100000;
    FSM_fft_64_stage_6_0_t652 = FSM_fft_64_stage_6_0_t651[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t653 = 32'b0;
    FSM_fft_64_stage_6_0_t654 = FSM_fft_64_stage_6_0_t653[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t655 = i_data_in_imag[FSM_fft_64_stage_6_0_t654 * 32 +: 32];
    FSM_fft_64_stage_6_0_t656 = 32'b00000000000000000000000000100000;
    FSM_fft_64_stage_6_0_t657 = FSM_fft_64_stage_6_0_t656[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t658 = i_data_in_imag[FSM_fft_64_stage_6_0_t657 * 32 +: 32];
    FSM_fft_64_stage_6_0_t659 = FSM_fft_64_stage_6_0_t650;
    FSM_fft_64_stage_6_0_t659[FSM_fft_64_stage_6_0_t652 * 32 +: 32] = FSM_fft_64_stage_6_0_t655 - FSM_fft_64_stage_6_0_t658;
    FSM_fft_64_stage_6_0_t660 = 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_6_0_t661 = FSM_fft_64_stage_6_0_t660[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t662 = 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_6_0_t663 = FSM_fft_64_stage_6_0_t662[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t664 = i_data_in_imag[FSM_fft_64_stage_6_0_t663 * 32 +: 32];
    FSM_fft_64_stage_6_0_t665 = 32'b00000000000000000000000000100001;
    FSM_fft_64_stage_6_0_t666 = FSM_fft_64_stage_6_0_t665[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t667 = i_data_in_imag[FSM_fft_64_stage_6_0_t666 * 32 +: 32];
    FSM_fft_64_stage_6_0_t668 = FSM_fft_64_stage_6_0_t664 + FSM_fft_64_stage_6_0_t667;
    FSM_fft_64_stage_6_0_t669 = FSM_fft_64_stage_6_0_t668[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t670 = FSM_fft_64_stage_6_0_t659;
    FSM_fft_64_stage_6_0_t670[FSM_fft_64_stage_6_0_t661 * 32 +: 32] = FSM_fft_64_stage_6_0_t669;
    FSM_fft_64_stage_6_0_t671 = 32'b00000000000000000000000000100001;
    FSM_fft_64_stage_6_0_t672 = FSM_fft_64_stage_6_0_t671[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t673 = 32'b00000000000000000000000000000001;
    FSM_fft_64_stage_6_0_t674 = FSM_fft_64_stage_6_0_t673[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t675 = i_data_in_imag[FSM_fft_64_stage_6_0_t674 * 32 +: 32];
    FSM_fft_64_stage_6_0_t676 = 32'b00000000000000000000000000100001;
    FSM_fft_64_stage_6_0_t677 = FSM_fft_64_stage_6_0_t676[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t678 = i_data_in_imag[FSM_fft_64_stage_6_0_t677 * 32 +: 32];
    FSM_fft_64_stage_6_0_t679 = FSM_fft_64_stage_6_0_t670;
    FSM_fft_64_stage_6_0_t679[FSM_fft_64_stage_6_0_t672 * 32 +: 32] = FSM_fft_64_stage_6_0_t675 - FSM_fft_64_stage_6_0_t678;
    FSM_fft_64_stage_6_0_t680 = 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_6_0_t681 = FSM_fft_64_stage_6_0_t680[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t682 = 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_6_0_t683 = FSM_fft_64_stage_6_0_t682[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t684 = i_data_in_imag[FSM_fft_64_stage_6_0_t683 * 32 +: 32];
    FSM_fft_64_stage_6_0_t685 = 32'b00000000000000000000000000100010;
    FSM_fft_64_stage_6_0_t686 = FSM_fft_64_stage_6_0_t685[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t687 = i_data_in_imag[FSM_fft_64_stage_6_0_t686 * 32 +: 32];
    FSM_fft_64_stage_6_0_t688 = FSM_fft_64_stage_6_0_t684 + FSM_fft_64_stage_6_0_t687;
    FSM_fft_64_stage_6_0_t689 = FSM_fft_64_stage_6_0_t688[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t690 = FSM_fft_64_stage_6_0_t679;
    FSM_fft_64_stage_6_0_t690[FSM_fft_64_stage_6_0_t681 * 32 +: 32] = FSM_fft_64_stage_6_0_t689;
    FSM_fft_64_stage_6_0_t691 = 32'b00000000000000000000000000100010;
    FSM_fft_64_stage_6_0_t692 = FSM_fft_64_stage_6_0_t691[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t693 = 32'b00000000000000000000000000000010;
    FSM_fft_64_stage_6_0_t694 = FSM_fft_64_stage_6_0_t693[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t695 = i_data_in_imag[FSM_fft_64_stage_6_0_t694 * 32 +: 32];
    FSM_fft_64_stage_6_0_t696 = 32'b00000000000000000000000000100010;
    FSM_fft_64_stage_6_0_t697 = FSM_fft_64_stage_6_0_t696[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t698 = i_data_in_imag[FSM_fft_64_stage_6_0_t697 * 32 +: 32];
    FSM_fft_64_stage_6_0_t699 = FSM_fft_64_stage_6_0_t690;
    FSM_fft_64_stage_6_0_t699[FSM_fft_64_stage_6_0_t692 * 32 +: 32] = FSM_fft_64_stage_6_0_t695 - FSM_fft_64_stage_6_0_t698;
    FSM_fft_64_stage_6_0_t700 = 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_6_0_t701 = FSM_fft_64_stage_6_0_t700[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t702 = 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_6_0_t703 = FSM_fft_64_stage_6_0_t702[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t704 = i_data_in_imag[FSM_fft_64_stage_6_0_t703 * 32 +: 32];
    FSM_fft_64_stage_6_0_t705 = 32'b00000000000000000000000000100011;
    FSM_fft_64_stage_6_0_t706 = FSM_fft_64_stage_6_0_t705[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t707 = i_data_in_imag[FSM_fft_64_stage_6_0_t706 * 32 +: 32];
    FSM_fft_64_stage_6_0_t708 = FSM_fft_64_stage_6_0_t704 + FSM_fft_64_stage_6_0_t707;
    FSM_fft_64_stage_6_0_t709 = FSM_fft_64_stage_6_0_t708[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t710 = FSM_fft_64_stage_6_0_t699;
    FSM_fft_64_stage_6_0_t710[FSM_fft_64_stage_6_0_t701 * 32 +: 32] = FSM_fft_64_stage_6_0_t709;
    FSM_fft_64_stage_6_0_t711 = 32'b00000000000000000000000000100011;
    FSM_fft_64_stage_6_0_t712 = FSM_fft_64_stage_6_0_t711[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t713 = 32'b00000000000000000000000000000011;
    FSM_fft_64_stage_6_0_t714 = FSM_fft_64_stage_6_0_t713[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t715 = i_data_in_imag[FSM_fft_64_stage_6_0_t714 * 32 +: 32];
    FSM_fft_64_stage_6_0_t716 = 32'b00000000000000000000000000100011;
    FSM_fft_64_stage_6_0_t717 = FSM_fft_64_stage_6_0_t716[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t718 = i_data_in_imag[FSM_fft_64_stage_6_0_t717 * 32 +: 32];
    FSM_fft_64_stage_6_0_t719 = FSM_fft_64_stage_6_0_t710;
    FSM_fft_64_stage_6_0_t719[FSM_fft_64_stage_6_0_t712 * 32 +: 32] = FSM_fft_64_stage_6_0_t715 - FSM_fft_64_stage_6_0_t718;
    FSM_fft_64_stage_6_0_t720 = 32'b00000000000000000000000000000100;
    FSM_fft_64_stage_6_0_t721 = FSM_fft_64_stage_6_0_t720[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t722 = 32'b00000000000000000000000000000100;
    FSM_fft_64_stage_6_0_t723 = FSM_fft_64_stage_6_0_t722[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t724 = i_data_in_imag[FSM_fft_64_stage_6_0_t723 * 32 +: 32];
    FSM_fft_64_stage_6_0_t725 = 32'b00000000000000000000000000100100;
    FSM_fft_64_stage_6_0_t726 = FSM_fft_64_stage_6_0_t725[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t727 = i_data_in_imag[FSM_fft_64_stage_6_0_t726 * 32 +: 32];
    FSM_fft_64_stage_6_0_t728 = FSM_fft_64_stage_6_0_t724 + FSM_fft_64_stage_6_0_t727;
    FSM_fft_64_stage_6_0_t729 = FSM_fft_64_stage_6_0_t728[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t730 = FSM_fft_64_stage_6_0_t719;
    FSM_fft_64_stage_6_0_t730[FSM_fft_64_stage_6_0_t721 * 32 +: 32] = FSM_fft_64_stage_6_0_t729;
    FSM_fft_64_stage_6_0_t731 = 32'b00000000000000000000000000100100;
    FSM_fft_64_stage_6_0_t732 = FSM_fft_64_stage_6_0_t731[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t733 = 32'b00000000000000000000000000000100;
    FSM_fft_64_stage_6_0_t734 = FSM_fft_64_stage_6_0_t733[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t735 = i_data_in_imag[FSM_fft_64_stage_6_0_t734 * 32 +: 32];
    FSM_fft_64_stage_6_0_t736 = 32'b00000000000000000000000000100100;
    FSM_fft_64_stage_6_0_t737 = FSM_fft_64_stage_6_0_t736[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t738 = i_data_in_imag[FSM_fft_64_stage_6_0_t737 * 32 +: 32];
    FSM_fft_64_stage_6_0_t739 = FSM_fft_64_stage_6_0_t730;
    FSM_fft_64_stage_6_0_t739[FSM_fft_64_stage_6_0_t732 * 32 +: 32] = FSM_fft_64_stage_6_0_t735 - FSM_fft_64_stage_6_0_t738;
    FSM_fft_64_stage_6_0_t740 = 32'b00000000000000000000000000000101;
    FSM_fft_64_stage_6_0_t741 = FSM_fft_64_stage_6_0_t740[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t742 = 32'b00000000000000000000000000000101;
    FSM_fft_64_stage_6_0_t743 = FSM_fft_64_stage_6_0_t742[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t744 = i_data_in_imag[FSM_fft_64_stage_6_0_t743 * 32 +: 32];
    FSM_fft_64_stage_6_0_t745 = 32'b00000000000000000000000000100101;
    FSM_fft_64_stage_6_0_t746 = FSM_fft_64_stage_6_0_t745[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t747 = i_data_in_imag[FSM_fft_64_stage_6_0_t746 * 32 +: 32];
    FSM_fft_64_stage_6_0_t748 = FSM_fft_64_stage_6_0_t744 + FSM_fft_64_stage_6_0_t747;
    FSM_fft_64_stage_6_0_t749 = FSM_fft_64_stage_6_0_t748[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t750 = FSM_fft_64_stage_6_0_t739;
    FSM_fft_64_stage_6_0_t750[FSM_fft_64_stage_6_0_t741 * 32 +: 32] = FSM_fft_64_stage_6_0_t749;
    FSM_fft_64_stage_6_0_t751 = 32'b00000000000000000000000000100101;
    FSM_fft_64_stage_6_0_t752 = FSM_fft_64_stage_6_0_t751[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t753 = 32'b00000000000000000000000000000101;
    FSM_fft_64_stage_6_0_t754 = FSM_fft_64_stage_6_0_t753[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t755 = i_data_in_imag[FSM_fft_64_stage_6_0_t754 * 32 +: 32];
    FSM_fft_64_stage_6_0_t756 = 32'b00000000000000000000000000100101;
    FSM_fft_64_stage_6_0_t757 = FSM_fft_64_stage_6_0_t756[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t758 = i_data_in_imag[FSM_fft_64_stage_6_0_t757 * 32 +: 32];
    FSM_fft_64_stage_6_0_t759 = FSM_fft_64_stage_6_0_t750;
    FSM_fft_64_stage_6_0_t759[FSM_fft_64_stage_6_0_t752 * 32 +: 32] = FSM_fft_64_stage_6_0_t755 - FSM_fft_64_stage_6_0_t758;
    FSM_fft_64_stage_6_0_t760 = 32'b00000000000000000000000000000110;
    FSM_fft_64_stage_6_0_t761 = FSM_fft_64_stage_6_0_t760[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t762 = 32'b00000000000000000000000000000110;
    FSM_fft_64_stage_6_0_t763 = FSM_fft_64_stage_6_0_t762[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t764 = i_data_in_imag[FSM_fft_64_stage_6_0_t763 * 32 +: 32];
    FSM_fft_64_stage_6_0_t765 = 32'b00000000000000000000000000100110;
    FSM_fft_64_stage_6_0_t766 = FSM_fft_64_stage_6_0_t765[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t767 = i_data_in_imag[FSM_fft_64_stage_6_0_t766 * 32 +: 32];
    FSM_fft_64_stage_6_0_t768 = FSM_fft_64_stage_6_0_t764 + FSM_fft_64_stage_6_0_t767;
    FSM_fft_64_stage_6_0_t769 = FSM_fft_64_stage_6_0_t768[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t770 = FSM_fft_64_stage_6_0_t759;
    FSM_fft_64_stage_6_0_t770[FSM_fft_64_stage_6_0_t761 * 32 +: 32] = FSM_fft_64_stage_6_0_t769;
    FSM_fft_64_stage_6_0_t771 = 32'b00000000000000000000000000100110;
    FSM_fft_64_stage_6_0_t772 = FSM_fft_64_stage_6_0_t771[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t773 = 32'b00000000000000000000000000000110;
    FSM_fft_64_stage_6_0_t774 = FSM_fft_64_stage_6_0_t773[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t775 = i_data_in_imag[FSM_fft_64_stage_6_0_t774 * 32 +: 32];
    FSM_fft_64_stage_6_0_t776 = 32'b00000000000000000000000000100110;
    FSM_fft_64_stage_6_0_t777 = FSM_fft_64_stage_6_0_t776[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t778 = i_data_in_imag[FSM_fft_64_stage_6_0_t777 * 32 +: 32];
    FSM_fft_64_stage_6_0_t779 = FSM_fft_64_stage_6_0_t770;
    FSM_fft_64_stage_6_0_t779[FSM_fft_64_stage_6_0_t772 * 32 +: 32] = FSM_fft_64_stage_6_0_t775 - FSM_fft_64_stage_6_0_t778;
    FSM_fft_64_stage_6_0_t780 = 32'b00000000000000000000000000000111;
    FSM_fft_64_stage_6_0_t781 = FSM_fft_64_stage_6_0_t780[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t782 = 32'b00000000000000000000000000000111;
    FSM_fft_64_stage_6_0_t783 = FSM_fft_64_stage_6_0_t782[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t784 = i_data_in_imag[FSM_fft_64_stage_6_0_t783 * 32 +: 32];
    FSM_fft_64_stage_6_0_t785 = 32'b00000000000000000000000000100111;
    FSM_fft_64_stage_6_0_t786 = FSM_fft_64_stage_6_0_t785[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t787 = i_data_in_imag[FSM_fft_64_stage_6_0_t786 * 32 +: 32];
    FSM_fft_64_stage_6_0_t788 = FSM_fft_64_stage_6_0_t784 + FSM_fft_64_stage_6_0_t787;
    FSM_fft_64_stage_6_0_t789 = FSM_fft_64_stage_6_0_t788[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t790 = FSM_fft_64_stage_6_0_t779;
    FSM_fft_64_stage_6_0_t790[FSM_fft_64_stage_6_0_t781 * 32 +: 32] = FSM_fft_64_stage_6_0_t789;
    FSM_fft_64_stage_6_0_t791 = 32'b00000000000000000000000000100111;
    FSM_fft_64_stage_6_0_t792 = FSM_fft_64_stage_6_0_t791[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t793 = 32'b00000000000000000000000000000111;
    FSM_fft_64_stage_6_0_t794 = FSM_fft_64_stage_6_0_t793[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t795 = i_data_in_imag[FSM_fft_64_stage_6_0_t794 * 32 +: 32];
    FSM_fft_64_stage_6_0_t796 = 32'b00000000000000000000000000100111;
    FSM_fft_64_stage_6_0_t797 = FSM_fft_64_stage_6_0_t796[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t798 = i_data_in_imag[FSM_fft_64_stage_6_0_t797 * 32 +: 32];
    FSM_fft_64_stage_6_0_t799 = FSM_fft_64_stage_6_0_t790;
    FSM_fft_64_stage_6_0_t799[FSM_fft_64_stage_6_0_t792 * 32 +: 32] = FSM_fft_64_stage_6_0_t795 - FSM_fft_64_stage_6_0_t798;
    FSM_fft_64_stage_6_0_t800 = 32'b00000000000000000000000000001000;
    FSM_fft_64_stage_6_0_t801 = FSM_fft_64_stage_6_0_t800[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t802 = 32'b00000000000000000000000000001000;
    FSM_fft_64_stage_6_0_t803 = FSM_fft_64_stage_6_0_t802[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t804 = i_data_in_imag[FSM_fft_64_stage_6_0_t803 * 32 +: 32];
    FSM_fft_64_stage_6_0_t805 = 32'b00000000000000000000000000101000;
    FSM_fft_64_stage_6_0_t806 = FSM_fft_64_stage_6_0_t805[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t807 = i_data_in_imag[FSM_fft_64_stage_6_0_t806 * 32 +: 32];
    FSM_fft_64_stage_6_0_t808 = FSM_fft_64_stage_6_0_t804 + FSM_fft_64_stage_6_0_t807;
    FSM_fft_64_stage_6_0_t809 = FSM_fft_64_stage_6_0_t808[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t810 = FSM_fft_64_stage_6_0_t799;
    FSM_fft_64_stage_6_0_t810[FSM_fft_64_stage_6_0_t801 * 32 +: 32] = FSM_fft_64_stage_6_0_t809;
    FSM_fft_64_stage_6_0_t811 = 32'b00000000000000000000000000101000;
    FSM_fft_64_stage_6_0_t812 = FSM_fft_64_stage_6_0_t811[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t813 = 32'b00000000000000000000000000001000;
    FSM_fft_64_stage_6_0_t814 = FSM_fft_64_stage_6_0_t813[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t815 = i_data_in_imag[FSM_fft_64_stage_6_0_t814 * 32 +: 32];
    FSM_fft_64_stage_6_0_t816 = 32'b00000000000000000000000000101000;
    FSM_fft_64_stage_6_0_t817 = FSM_fft_64_stage_6_0_t816[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t818 = i_data_in_imag[FSM_fft_64_stage_6_0_t817 * 32 +: 32];
    FSM_fft_64_stage_6_0_t819 = FSM_fft_64_stage_6_0_t810;
    FSM_fft_64_stage_6_0_t819[FSM_fft_64_stage_6_0_t812 * 32 +: 32] = FSM_fft_64_stage_6_0_t815 - FSM_fft_64_stage_6_0_t818;
    FSM_fft_64_stage_6_0_t820 = 32'b00000000000000000000000000001001;
    FSM_fft_64_stage_6_0_t821 = FSM_fft_64_stage_6_0_t820[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t822 = 32'b00000000000000000000000000001001;
    FSM_fft_64_stage_6_0_t823 = FSM_fft_64_stage_6_0_t822[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t824 = i_data_in_imag[FSM_fft_64_stage_6_0_t823 * 32 +: 32];
    FSM_fft_64_stage_6_0_t825 = 32'b00000000000000000000000000101001;
    FSM_fft_64_stage_6_0_t826 = FSM_fft_64_stage_6_0_t825[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t827 = i_data_in_imag[FSM_fft_64_stage_6_0_t826 * 32 +: 32];
    FSM_fft_64_stage_6_0_t828 = FSM_fft_64_stage_6_0_t824 + FSM_fft_64_stage_6_0_t827;
    FSM_fft_64_stage_6_0_t829 = FSM_fft_64_stage_6_0_t828[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t830 = FSM_fft_64_stage_6_0_t819;
    FSM_fft_64_stage_6_0_t830[FSM_fft_64_stage_6_0_t821 * 32 +: 32] = FSM_fft_64_stage_6_0_t829;
    FSM_fft_64_stage_6_0_t831 = 32'b00000000000000000000000000101001;
    FSM_fft_64_stage_6_0_t832 = FSM_fft_64_stage_6_0_t831[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t833 = 32'b00000000000000000000000000001001;
    FSM_fft_64_stage_6_0_t834 = FSM_fft_64_stage_6_0_t833[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t835 = i_data_in_imag[FSM_fft_64_stage_6_0_t834 * 32 +: 32];
    FSM_fft_64_stage_6_0_t836 = 32'b00000000000000000000000000101001;
    FSM_fft_64_stage_6_0_t837 = FSM_fft_64_stage_6_0_t836[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t838 = i_data_in_imag[FSM_fft_64_stage_6_0_t837 * 32 +: 32];
    FSM_fft_64_stage_6_0_t839 = FSM_fft_64_stage_6_0_t830;
    FSM_fft_64_stage_6_0_t839[FSM_fft_64_stage_6_0_t832 * 32 +: 32] = FSM_fft_64_stage_6_0_t835 - FSM_fft_64_stage_6_0_t838;
    FSM_fft_64_stage_6_0_t840 = 32'b00000000000000000000000000001010;
    FSM_fft_64_stage_6_0_t841 = FSM_fft_64_stage_6_0_t840[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t842 = 32'b00000000000000000000000000001010;
    FSM_fft_64_stage_6_0_t843 = FSM_fft_64_stage_6_0_t842[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t844 = i_data_in_imag[FSM_fft_64_stage_6_0_t843 * 32 +: 32];
    FSM_fft_64_stage_6_0_t845 = 32'b00000000000000000000000000101010;
    FSM_fft_64_stage_6_0_t846 = FSM_fft_64_stage_6_0_t845[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t847 = i_data_in_imag[FSM_fft_64_stage_6_0_t846 * 32 +: 32];
    FSM_fft_64_stage_6_0_t848 = FSM_fft_64_stage_6_0_t844 + FSM_fft_64_stage_6_0_t847;
    FSM_fft_64_stage_6_0_t849 = FSM_fft_64_stage_6_0_t848[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t850 = FSM_fft_64_stage_6_0_t839;
    FSM_fft_64_stage_6_0_t850[FSM_fft_64_stage_6_0_t841 * 32 +: 32] = FSM_fft_64_stage_6_0_t849;
    FSM_fft_64_stage_6_0_t851 = 32'b00000000000000000000000000101010;
    FSM_fft_64_stage_6_0_t852 = FSM_fft_64_stage_6_0_t851[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t853 = 32'b00000000000000000000000000001010;
    FSM_fft_64_stage_6_0_t854 = FSM_fft_64_stage_6_0_t853[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t855 = i_data_in_imag[FSM_fft_64_stage_6_0_t854 * 32 +: 32];
    FSM_fft_64_stage_6_0_t856 = 32'b00000000000000000000000000101010;
    FSM_fft_64_stage_6_0_t857 = FSM_fft_64_stage_6_0_t856[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t858 = i_data_in_imag[FSM_fft_64_stage_6_0_t857 * 32 +: 32];
    FSM_fft_64_stage_6_0_t859 = FSM_fft_64_stage_6_0_t850;
    FSM_fft_64_stage_6_0_t859[FSM_fft_64_stage_6_0_t852 * 32 +: 32] = FSM_fft_64_stage_6_0_t855 - FSM_fft_64_stage_6_0_t858;
    FSM_fft_64_stage_6_0_t860 = 32'b00000000000000000000000000001011;
    FSM_fft_64_stage_6_0_t861 = FSM_fft_64_stage_6_0_t860[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t862 = 32'b00000000000000000000000000001011;
    FSM_fft_64_stage_6_0_t863 = FSM_fft_64_stage_6_0_t862[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t864 = i_data_in_imag[FSM_fft_64_stage_6_0_t863 * 32 +: 32];
    FSM_fft_64_stage_6_0_t865 = 32'b00000000000000000000000000101011;
    FSM_fft_64_stage_6_0_t866 = FSM_fft_64_stage_6_0_t865[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t867 = i_data_in_imag[FSM_fft_64_stage_6_0_t866 * 32 +: 32];
    FSM_fft_64_stage_6_0_t868 = FSM_fft_64_stage_6_0_t864 + FSM_fft_64_stage_6_0_t867;
    FSM_fft_64_stage_6_0_t869 = FSM_fft_64_stage_6_0_t868[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t870 = FSM_fft_64_stage_6_0_t859;
    FSM_fft_64_stage_6_0_t870[FSM_fft_64_stage_6_0_t861 * 32 +: 32] = FSM_fft_64_stage_6_0_t869;
    FSM_fft_64_stage_6_0_t871 = 32'b00000000000000000000000000101011;
    FSM_fft_64_stage_6_0_t872 = FSM_fft_64_stage_6_0_t871[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t873 = 32'b00000000000000000000000000001011;
    FSM_fft_64_stage_6_0_t874 = FSM_fft_64_stage_6_0_t873[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t875 = i_data_in_imag[FSM_fft_64_stage_6_0_t874 * 32 +: 32];
    FSM_fft_64_stage_6_0_t876 = 32'b00000000000000000000000000101011;
    FSM_fft_64_stage_6_0_t877 = FSM_fft_64_stage_6_0_t876[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t878 = i_data_in_imag[FSM_fft_64_stage_6_0_t877 * 32 +: 32];
    FSM_fft_64_stage_6_0_t879 = FSM_fft_64_stage_6_0_t870;
    FSM_fft_64_stage_6_0_t879[FSM_fft_64_stage_6_0_t872 * 32 +: 32] = FSM_fft_64_stage_6_0_t875 - FSM_fft_64_stage_6_0_t878;
    FSM_fft_64_stage_6_0_t880 = 32'b00000000000000000000000000001100;
    FSM_fft_64_stage_6_0_t881 = FSM_fft_64_stage_6_0_t880[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t882 = 32'b00000000000000000000000000001100;
    FSM_fft_64_stage_6_0_t883 = FSM_fft_64_stage_6_0_t882[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t884 = i_data_in_imag[FSM_fft_64_stage_6_0_t883 * 32 +: 32];
    FSM_fft_64_stage_6_0_t885 = 32'b00000000000000000000000000101100;
    FSM_fft_64_stage_6_0_t886 = FSM_fft_64_stage_6_0_t885[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t887 = i_data_in_imag[FSM_fft_64_stage_6_0_t886 * 32 +: 32];
    FSM_fft_64_stage_6_0_t888 = FSM_fft_64_stage_6_0_t884 + FSM_fft_64_stage_6_0_t887;
    FSM_fft_64_stage_6_0_t889 = FSM_fft_64_stage_6_0_t888[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t890 = FSM_fft_64_stage_6_0_t879;
    FSM_fft_64_stage_6_0_t890[FSM_fft_64_stage_6_0_t881 * 32 +: 32] = FSM_fft_64_stage_6_0_t889;
    FSM_fft_64_stage_6_0_t891 = 32'b00000000000000000000000000101100;
    FSM_fft_64_stage_6_0_t892 = FSM_fft_64_stage_6_0_t891[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t893 = 32'b00000000000000000000000000001100;
    FSM_fft_64_stage_6_0_t894 = FSM_fft_64_stage_6_0_t893[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t895 = i_data_in_imag[FSM_fft_64_stage_6_0_t894 * 32 +: 32];
    FSM_fft_64_stage_6_0_t896 = 32'b00000000000000000000000000101100;
    FSM_fft_64_stage_6_0_t897 = FSM_fft_64_stage_6_0_t896[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t898 = i_data_in_imag[FSM_fft_64_stage_6_0_t897 * 32 +: 32];
    FSM_fft_64_stage_6_0_t899 = FSM_fft_64_stage_6_0_t890;
    FSM_fft_64_stage_6_0_t899[FSM_fft_64_stage_6_0_t892 * 32 +: 32] = FSM_fft_64_stage_6_0_t895 - FSM_fft_64_stage_6_0_t898;
    FSM_fft_64_stage_6_0_t900 = 32'b00000000000000000000000000001101;
    FSM_fft_64_stage_6_0_t901 = FSM_fft_64_stage_6_0_t900[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t902 = 32'b00000000000000000000000000001101;
    FSM_fft_64_stage_6_0_t903 = FSM_fft_64_stage_6_0_t902[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t904 = i_data_in_imag[FSM_fft_64_stage_6_0_t903 * 32 +: 32];
    FSM_fft_64_stage_6_0_t905 = 32'b00000000000000000000000000101101;
    FSM_fft_64_stage_6_0_t906 = FSM_fft_64_stage_6_0_t905[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t907 = i_data_in_imag[FSM_fft_64_stage_6_0_t906 * 32 +: 32];
    FSM_fft_64_stage_6_0_t908 = FSM_fft_64_stage_6_0_t904 + FSM_fft_64_stage_6_0_t907;
    FSM_fft_64_stage_6_0_t909 = FSM_fft_64_stage_6_0_t908[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t910 = FSM_fft_64_stage_6_0_t899;
    FSM_fft_64_stage_6_0_t910[FSM_fft_64_stage_6_0_t901 * 32 +: 32] = FSM_fft_64_stage_6_0_t909;
    FSM_fft_64_stage_6_0_t911 = 32'b00000000000000000000000000101101;
    FSM_fft_64_stage_6_0_t912 = FSM_fft_64_stage_6_0_t911[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t913 = 32'b00000000000000000000000000001101;
    FSM_fft_64_stage_6_0_t914 = FSM_fft_64_stage_6_0_t913[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t915 = i_data_in_imag[FSM_fft_64_stage_6_0_t914 * 32 +: 32];
    FSM_fft_64_stage_6_0_t916 = 32'b00000000000000000000000000101101;
    FSM_fft_64_stage_6_0_t917 = FSM_fft_64_stage_6_0_t916[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t918 = i_data_in_imag[FSM_fft_64_stage_6_0_t917 * 32 +: 32];
    FSM_fft_64_stage_6_0_t919 = FSM_fft_64_stage_6_0_t910;
    FSM_fft_64_stage_6_0_t919[FSM_fft_64_stage_6_0_t912 * 32 +: 32] = FSM_fft_64_stage_6_0_t915 - FSM_fft_64_stage_6_0_t918;
    FSM_fft_64_stage_6_0_t920 = 32'b00000000000000000000000000001110;
    FSM_fft_64_stage_6_0_t921 = FSM_fft_64_stage_6_0_t920[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t922 = 32'b00000000000000000000000000001110;
    FSM_fft_64_stage_6_0_t923 = FSM_fft_64_stage_6_0_t922[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t924 = i_data_in_imag[FSM_fft_64_stage_6_0_t923 * 32 +: 32];
    FSM_fft_64_stage_6_0_t925 = 32'b00000000000000000000000000101110;
    FSM_fft_64_stage_6_0_t926 = FSM_fft_64_stage_6_0_t925[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t927 = i_data_in_imag[FSM_fft_64_stage_6_0_t926 * 32 +: 32];
    FSM_fft_64_stage_6_0_t928 = FSM_fft_64_stage_6_0_t924 + FSM_fft_64_stage_6_0_t927;
    FSM_fft_64_stage_6_0_t929 = FSM_fft_64_stage_6_0_t928[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t930 = FSM_fft_64_stage_6_0_t919;
    FSM_fft_64_stage_6_0_t930[FSM_fft_64_stage_6_0_t921 * 32 +: 32] = FSM_fft_64_stage_6_0_t929;
    FSM_fft_64_stage_6_0_t931 = 32'b00000000000000000000000000101110;
    FSM_fft_64_stage_6_0_t932 = FSM_fft_64_stage_6_0_t931[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t933 = 32'b00000000000000000000000000001110;
    FSM_fft_64_stage_6_0_t934 = FSM_fft_64_stage_6_0_t933[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t935 = i_data_in_imag[FSM_fft_64_stage_6_0_t934 * 32 +: 32];
    FSM_fft_64_stage_6_0_t936 = 32'b00000000000000000000000000101110;
    FSM_fft_64_stage_6_0_t937 = FSM_fft_64_stage_6_0_t936[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t938 = i_data_in_imag[FSM_fft_64_stage_6_0_t937 * 32 +: 32];
    FSM_fft_64_stage_6_0_t939 = FSM_fft_64_stage_6_0_t930;
    FSM_fft_64_stage_6_0_t939[FSM_fft_64_stage_6_0_t932 * 32 +: 32] = FSM_fft_64_stage_6_0_t935 - FSM_fft_64_stage_6_0_t938;
    FSM_fft_64_stage_6_0_t940 = 32'b00000000000000000000000000001111;
    FSM_fft_64_stage_6_0_t941 = FSM_fft_64_stage_6_0_t940[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t942 = 32'b00000000000000000000000000001111;
    FSM_fft_64_stage_6_0_t943 = FSM_fft_64_stage_6_0_t942[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t944 = i_data_in_imag[FSM_fft_64_stage_6_0_t943 * 32 +: 32];
    FSM_fft_64_stage_6_0_t945 = 32'b00000000000000000000000000101111;
    FSM_fft_64_stage_6_0_t946 = FSM_fft_64_stage_6_0_t945[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t947 = i_data_in_imag[FSM_fft_64_stage_6_0_t946 * 32 +: 32];
    FSM_fft_64_stage_6_0_t948 = FSM_fft_64_stage_6_0_t944 + FSM_fft_64_stage_6_0_t947;
    FSM_fft_64_stage_6_0_t949 = FSM_fft_64_stage_6_0_t948[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t950 = FSM_fft_64_stage_6_0_t939;
    FSM_fft_64_stage_6_0_t950[FSM_fft_64_stage_6_0_t941 * 32 +: 32] = FSM_fft_64_stage_6_0_t949;
    FSM_fft_64_stage_6_0_t951 = 32'b00000000000000000000000000101111;
    FSM_fft_64_stage_6_0_t952 = FSM_fft_64_stage_6_0_t951[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t953 = 32'b00000000000000000000000000001111;
    FSM_fft_64_stage_6_0_t954 = FSM_fft_64_stage_6_0_t953[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t955 = i_data_in_imag[FSM_fft_64_stage_6_0_t954 * 32 +: 32];
    FSM_fft_64_stage_6_0_t956 = 32'b00000000000000000000000000101111;
    FSM_fft_64_stage_6_0_t957 = FSM_fft_64_stage_6_0_t956[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t958 = i_data_in_imag[FSM_fft_64_stage_6_0_t957 * 32 +: 32];
    FSM_fft_64_stage_6_0_t959 = FSM_fft_64_stage_6_0_t950;
    FSM_fft_64_stage_6_0_t959[FSM_fft_64_stage_6_0_t952 * 32 +: 32] = FSM_fft_64_stage_6_0_t955 - FSM_fft_64_stage_6_0_t958;
    FSM_fft_64_stage_6_0_t960 = 32'b00000000000000000000000000010000;
    FSM_fft_64_stage_6_0_t961 = FSM_fft_64_stage_6_0_t960[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t962 = 32'b00000000000000000000000000010000;
    FSM_fft_64_stage_6_0_t963 = FSM_fft_64_stage_6_0_t962[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t964 = i_data_in_imag[FSM_fft_64_stage_6_0_t963 * 32 +: 32];
    FSM_fft_64_stage_6_0_t965 = 32'b00000000000000000000000000110000;
    FSM_fft_64_stage_6_0_t966 = FSM_fft_64_stage_6_0_t965[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t967 = i_data_in_imag[FSM_fft_64_stage_6_0_t966 * 32 +: 32];
    FSM_fft_64_stage_6_0_t968 = FSM_fft_64_stage_6_0_t964 + FSM_fft_64_stage_6_0_t967;
    FSM_fft_64_stage_6_0_t969 = FSM_fft_64_stage_6_0_t968[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t970 = FSM_fft_64_stage_6_0_t959;
    FSM_fft_64_stage_6_0_t970[FSM_fft_64_stage_6_0_t961 * 32 +: 32] = FSM_fft_64_stage_6_0_t969;
    FSM_fft_64_stage_6_0_t971 = 32'b00000000000000000000000000110000;
    FSM_fft_64_stage_6_0_t972 = FSM_fft_64_stage_6_0_t971[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t973 = 32'b00000000000000000000000000010000;
    FSM_fft_64_stage_6_0_t974 = FSM_fft_64_stage_6_0_t973[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t975 = i_data_in_imag[FSM_fft_64_stage_6_0_t974 * 32 +: 32];
    FSM_fft_64_stage_6_0_t976 = 32'b00000000000000000000000000110000;
    FSM_fft_64_stage_6_0_t977 = FSM_fft_64_stage_6_0_t976[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t978 = i_data_in_imag[FSM_fft_64_stage_6_0_t977 * 32 +: 32];
    FSM_fft_64_stage_6_0_t979 = FSM_fft_64_stage_6_0_t970;
    FSM_fft_64_stage_6_0_t979[FSM_fft_64_stage_6_0_t972 * 32 +: 32] = FSM_fft_64_stage_6_0_t975 - FSM_fft_64_stage_6_0_t978;
    FSM_fft_64_stage_6_0_t980 = 32'b00000000000000000000000000010001;
    FSM_fft_64_stage_6_0_t981 = FSM_fft_64_stage_6_0_t980[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t982 = 32'b00000000000000000000000000010001;
    FSM_fft_64_stage_6_0_t983 = FSM_fft_64_stage_6_0_t982[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t984 = i_data_in_imag[FSM_fft_64_stage_6_0_t983 * 32 +: 32];
    FSM_fft_64_stage_6_0_t985 = 32'b00000000000000000000000000110001;
    FSM_fft_64_stage_6_0_t986 = FSM_fft_64_stage_6_0_t985[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t987 = i_data_in_imag[FSM_fft_64_stage_6_0_t986 * 32 +: 32];
    FSM_fft_64_stage_6_0_t988 = FSM_fft_64_stage_6_0_t984 + FSM_fft_64_stage_6_0_t987;
    FSM_fft_64_stage_6_0_t989 = FSM_fft_64_stage_6_0_t988[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t990 = FSM_fft_64_stage_6_0_t979;
    FSM_fft_64_stage_6_0_t990[FSM_fft_64_stage_6_0_t981 * 32 +: 32] = FSM_fft_64_stage_6_0_t989;
    FSM_fft_64_stage_6_0_t991 = 32'b00000000000000000000000000110001;
    FSM_fft_64_stage_6_0_t992 = FSM_fft_64_stage_6_0_t991[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t993 = 32'b00000000000000000000000000010001;
    FSM_fft_64_stage_6_0_t994 = FSM_fft_64_stage_6_0_t993[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t995 = i_data_in_imag[FSM_fft_64_stage_6_0_t994 * 32 +: 32];
    FSM_fft_64_stage_6_0_t996 = 32'b00000000000000000000000000110001;
    FSM_fft_64_stage_6_0_t997 = FSM_fft_64_stage_6_0_t996[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t998 = i_data_in_imag[FSM_fft_64_stage_6_0_t997 * 32 +: 32];
    FSM_fft_64_stage_6_0_t999 = FSM_fft_64_stage_6_0_t990;
    FSM_fft_64_stage_6_0_t999[FSM_fft_64_stage_6_0_t992 * 32 +: 32] = FSM_fft_64_stage_6_0_t995 - FSM_fft_64_stage_6_0_t998;
    FSM_fft_64_stage_6_0_t1000 = 32'b00000000000000000000000000010010;
    FSM_fft_64_stage_6_0_t1001 = FSM_fft_64_stage_6_0_t1000[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1002 = 32'b00000000000000000000000000010010;
    FSM_fft_64_stage_6_0_t1003 = FSM_fft_64_stage_6_0_t1002[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1004 = i_data_in_imag[FSM_fft_64_stage_6_0_t1003 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1005 = 32'b00000000000000000000000000110010;
    FSM_fft_64_stage_6_0_t1006 = FSM_fft_64_stage_6_0_t1005[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1007 = i_data_in_imag[FSM_fft_64_stage_6_0_t1006 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1008 = FSM_fft_64_stage_6_0_t1004 + FSM_fft_64_stage_6_0_t1007;
    FSM_fft_64_stage_6_0_t1009 = FSM_fft_64_stage_6_0_t1008[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t1010 = FSM_fft_64_stage_6_0_t999;
    FSM_fft_64_stage_6_0_t1010[FSM_fft_64_stage_6_0_t1001 * 32 +: 32] = FSM_fft_64_stage_6_0_t1009;
    FSM_fft_64_stage_6_0_t1011 = 32'b00000000000000000000000000110010;
    FSM_fft_64_stage_6_0_t1012 = FSM_fft_64_stage_6_0_t1011[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1013 = 32'b00000000000000000000000000010010;
    FSM_fft_64_stage_6_0_t1014 = FSM_fft_64_stage_6_0_t1013[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1015 = i_data_in_imag[FSM_fft_64_stage_6_0_t1014 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1016 = 32'b00000000000000000000000000110010;
    FSM_fft_64_stage_6_0_t1017 = FSM_fft_64_stage_6_0_t1016[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1018 = i_data_in_imag[FSM_fft_64_stage_6_0_t1017 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1019 = FSM_fft_64_stage_6_0_t1010;
    FSM_fft_64_stage_6_0_t1019[FSM_fft_64_stage_6_0_t1012 * 32 +: 32] = FSM_fft_64_stage_6_0_t1015 - FSM_fft_64_stage_6_0_t1018;
    FSM_fft_64_stage_6_0_t1020 = 32'b00000000000000000000000000010011;
    FSM_fft_64_stage_6_0_t1021 = FSM_fft_64_stage_6_0_t1020[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1022 = 32'b00000000000000000000000000010011;
    FSM_fft_64_stage_6_0_t1023 = FSM_fft_64_stage_6_0_t1022[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1024 = i_data_in_imag[FSM_fft_64_stage_6_0_t1023 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1025 = 32'b00000000000000000000000000110011;
    FSM_fft_64_stage_6_0_t1026 = FSM_fft_64_stage_6_0_t1025[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1027 = i_data_in_imag[FSM_fft_64_stage_6_0_t1026 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1028 = FSM_fft_64_stage_6_0_t1024 + FSM_fft_64_stage_6_0_t1027;
    FSM_fft_64_stage_6_0_t1029 = FSM_fft_64_stage_6_0_t1028[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t1030 = FSM_fft_64_stage_6_0_t1019;
    FSM_fft_64_stage_6_0_t1030[FSM_fft_64_stage_6_0_t1021 * 32 +: 32] = FSM_fft_64_stage_6_0_t1029;
    FSM_fft_64_stage_6_0_t1031 = 32'b00000000000000000000000000110011;
    FSM_fft_64_stage_6_0_t1032 = FSM_fft_64_stage_6_0_t1031[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1033 = 32'b00000000000000000000000000010011;
    FSM_fft_64_stage_6_0_t1034 = FSM_fft_64_stage_6_0_t1033[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1035 = i_data_in_imag[FSM_fft_64_stage_6_0_t1034 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1036 = 32'b00000000000000000000000000110011;
    FSM_fft_64_stage_6_0_t1037 = FSM_fft_64_stage_6_0_t1036[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1038 = i_data_in_imag[FSM_fft_64_stage_6_0_t1037 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1039 = FSM_fft_64_stage_6_0_t1030;
    FSM_fft_64_stage_6_0_t1039[FSM_fft_64_stage_6_0_t1032 * 32 +: 32] = FSM_fft_64_stage_6_0_t1035 - FSM_fft_64_stage_6_0_t1038;
    FSM_fft_64_stage_6_0_t1040 = 32'b00000000000000000000000000010100;
    FSM_fft_64_stage_6_0_t1041 = FSM_fft_64_stage_6_0_t1040[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1042 = 32'b00000000000000000000000000010100;
    FSM_fft_64_stage_6_0_t1043 = FSM_fft_64_stage_6_0_t1042[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1044 = i_data_in_imag[FSM_fft_64_stage_6_0_t1043 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1045 = 32'b00000000000000000000000000110100;
    FSM_fft_64_stage_6_0_t1046 = FSM_fft_64_stage_6_0_t1045[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1047 = i_data_in_imag[FSM_fft_64_stage_6_0_t1046 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1048 = FSM_fft_64_stage_6_0_t1044 + FSM_fft_64_stage_6_0_t1047;
    FSM_fft_64_stage_6_0_t1049 = FSM_fft_64_stage_6_0_t1048[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t1050 = FSM_fft_64_stage_6_0_t1039;
    FSM_fft_64_stage_6_0_t1050[FSM_fft_64_stage_6_0_t1041 * 32 +: 32] = FSM_fft_64_stage_6_0_t1049;
    FSM_fft_64_stage_6_0_t1051 = 32'b00000000000000000000000000110100;
    FSM_fft_64_stage_6_0_t1052 = FSM_fft_64_stage_6_0_t1051[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1053 = 32'b00000000000000000000000000010100;
    FSM_fft_64_stage_6_0_t1054 = FSM_fft_64_stage_6_0_t1053[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1055 = i_data_in_imag[FSM_fft_64_stage_6_0_t1054 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1056 = 32'b00000000000000000000000000110100;
    FSM_fft_64_stage_6_0_t1057 = FSM_fft_64_stage_6_0_t1056[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1058 = i_data_in_imag[FSM_fft_64_stage_6_0_t1057 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1059 = FSM_fft_64_stage_6_0_t1050;
    FSM_fft_64_stage_6_0_t1059[FSM_fft_64_stage_6_0_t1052 * 32 +: 32] = FSM_fft_64_stage_6_0_t1055 - FSM_fft_64_stage_6_0_t1058;
    FSM_fft_64_stage_6_0_t1060 = 32'b00000000000000000000000000010101;
    FSM_fft_64_stage_6_0_t1061 = FSM_fft_64_stage_6_0_t1060[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1062 = 32'b00000000000000000000000000010101;
    FSM_fft_64_stage_6_0_t1063 = FSM_fft_64_stage_6_0_t1062[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1064 = i_data_in_imag[FSM_fft_64_stage_6_0_t1063 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1065 = 32'b00000000000000000000000000110101;
    FSM_fft_64_stage_6_0_t1066 = FSM_fft_64_stage_6_0_t1065[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1067 = i_data_in_imag[FSM_fft_64_stage_6_0_t1066 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1068 = FSM_fft_64_stage_6_0_t1064 + FSM_fft_64_stage_6_0_t1067;
    FSM_fft_64_stage_6_0_t1069 = FSM_fft_64_stage_6_0_t1068[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t1070 = FSM_fft_64_stage_6_0_t1059;
    FSM_fft_64_stage_6_0_t1070[FSM_fft_64_stage_6_0_t1061 * 32 +: 32] = FSM_fft_64_stage_6_0_t1069;
    FSM_fft_64_stage_6_0_t1071 = 32'b00000000000000000000000000110101;
    FSM_fft_64_stage_6_0_t1072 = FSM_fft_64_stage_6_0_t1071[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1073 = 32'b00000000000000000000000000010101;
    FSM_fft_64_stage_6_0_t1074 = FSM_fft_64_stage_6_0_t1073[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1075 = i_data_in_imag[FSM_fft_64_stage_6_0_t1074 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1076 = 32'b00000000000000000000000000110101;
    FSM_fft_64_stage_6_0_t1077 = FSM_fft_64_stage_6_0_t1076[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1078 = i_data_in_imag[FSM_fft_64_stage_6_0_t1077 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1079 = FSM_fft_64_stage_6_0_t1070;
    FSM_fft_64_stage_6_0_t1079[FSM_fft_64_stage_6_0_t1072 * 32 +: 32] = FSM_fft_64_stage_6_0_t1075 - FSM_fft_64_stage_6_0_t1078;
    FSM_fft_64_stage_6_0_t1080 = 32'b00000000000000000000000000010110;
    FSM_fft_64_stage_6_0_t1081 = FSM_fft_64_stage_6_0_t1080[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1082 = 32'b00000000000000000000000000010110;
    FSM_fft_64_stage_6_0_t1083 = FSM_fft_64_stage_6_0_t1082[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1084 = i_data_in_imag[FSM_fft_64_stage_6_0_t1083 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1085 = 32'b00000000000000000000000000110110;
    FSM_fft_64_stage_6_0_t1086 = FSM_fft_64_stage_6_0_t1085[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1087 = i_data_in_imag[FSM_fft_64_stage_6_0_t1086 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1088 = FSM_fft_64_stage_6_0_t1084 + FSM_fft_64_stage_6_0_t1087;
    FSM_fft_64_stage_6_0_t1089 = FSM_fft_64_stage_6_0_t1088[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t1090 = FSM_fft_64_stage_6_0_t1079;
    FSM_fft_64_stage_6_0_t1090[FSM_fft_64_stage_6_0_t1081 * 32 +: 32] = FSM_fft_64_stage_6_0_t1089;
    FSM_fft_64_stage_6_0_t1091 = 32'b00000000000000000000000000110110;
    FSM_fft_64_stage_6_0_t1092 = FSM_fft_64_stage_6_0_t1091[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1093 = 32'b00000000000000000000000000010110;
    FSM_fft_64_stage_6_0_t1094 = FSM_fft_64_stage_6_0_t1093[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1095 = i_data_in_imag[FSM_fft_64_stage_6_0_t1094 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1096 = 32'b00000000000000000000000000110110;
    FSM_fft_64_stage_6_0_t1097 = FSM_fft_64_stage_6_0_t1096[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1098 = i_data_in_imag[FSM_fft_64_stage_6_0_t1097 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1099 = FSM_fft_64_stage_6_0_t1090;
    FSM_fft_64_stage_6_0_t1099[FSM_fft_64_stage_6_0_t1092 * 32 +: 32] = FSM_fft_64_stage_6_0_t1095 - FSM_fft_64_stage_6_0_t1098;
    FSM_fft_64_stage_6_0_t1100 = 32'b00000000000000000000000000010111;
    FSM_fft_64_stage_6_0_t1101 = FSM_fft_64_stage_6_0_t1100[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1102 = 32'b00000000000000000000000000010111;
    FSM_fft_64_stage_6_0_t1103 = FSM_fft_64_stage_6_0_t1102[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1104 = i_data_in_imag[FSM_fft_64_stage_6_0_t1103 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1105 = 32'b00000000000000000000000000110111;
    FSM_fft_64_stage_6_0_t1106 = FSM_fft_64_stage_6_0_t1105[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1107 = i_data_in_imag[FSM_fft_64_stage_6_0_t1106 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1108 = FSM_fft_64_stage_6_0_t1104 + FSM_fft_64_stage_6_0_t1107;
    FSM_fft_64_stage_6_0_t1109 = FSM_fft_64_stage_6_0_t1108[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t1110 = FSM_fft_64_stage_6_0_t1099;
    FSM_fft_64_stage_6_0_t1110[FSM_fft_64_stage_6_0_t1101 * 32 +: 32] = FSM_fft_64_stage_6_0_t1109;
    FSM_fft_64_stage_6_0_t1111 = 32'b00000000000000000000000000110111;
    FSM_fft_64_stage_6_0_t1112 = FSM_fft_64_stage_6_0_t1111[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1113 = 32'b00000000000000000000000000010111;
    FSM_fft_64_stage_6_0_t1114 = FSM_fft_64_stage_6_0_t1113[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1115 = i_data_in_imag[FSM_fft_64_stage_6_0_t1114 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1116 = 32'b00000000000000000000000000110111;
    FSM_fft_64_stage_6_0_t1117 = FSM_fft_64_stage_6_0_t1116[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1118 = i_data_in_imag[FSM_fft_64_stage_6_0_t1117 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1119 = FSM_fft_64_stage_6_0_t1110;
    FSM_fft_64_stage_6_0_t1119[FSM_fft_64_stage_6_0_t1112 * 32 +: 32] = FSM_fft_64_stage_6_0_t1115 - FSM_fft_64_stage_6_0_t1118;
    FSM_fft_64_stage_6_0_t1120 = 32'b00000000000000000000000000011000;
    FSM_fft_64_stage_6_0_t1121 = FSM_fft_64_stage_6_0_t1120[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1122 = 32'b00000000000000000000000000011000;
    FSM_fft_64_stage_6_0_t1123 = FSM_fft_64_stage_6_0_t1122[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1124 = i_data_in_imag[FSM_fft_64_stage_6_0_t1123 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1125 = 32'b00000000000000000000000000111000;
    FSM_fft_64_stage_6_0_t1126 = FSM_fft_64_stage_6_0_t1125[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1127 = i_data_in_imag[FSM_fft_64_stage_6_0_t1126 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1128 = FSM_fft_64_stage_6_0_t1124 + FSM_fft_64_stage_6_0_t1127;
    FSM_fft_64_stage_6_0_t1129 = FSM_fft_64_stage_6_0_t1128[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t1130 = FSM_fft_64_stage_6_0_t1119;
    FSM_fft_64_stage_6_0_t1130[FSM_fft_64_stage_6_0_t1121 * 32 +: 32] = FSM_fft_64_stage_6_0_t1129;
    FSM_fft_64_stage_6_0_t1131 = 32'b00000000000000000000000000111000;
    FSM_fft_64_stage_6_0_t1132 = FSM_fft_64_stage_6_0_t1131[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1133 = 32'b00000000000000000000000000011000;
    FSM_fft_64_stage_6_0_t1134 = FSM_fft_64_stage_6_0_t1133[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1135 = i_data_in_imag[FSM_fft_64_stage_6_0_t1134 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1136 = 32'b00000000000000000000000000111000;
    FSM_fft_64_stage_6_0_t1137 = FSM_fft_64_stage_6_0_t1136[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1138 = i_data_in_imag[FSM_fft_64_stage_6_0_t1137 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1139 = FSM_fft_64_stage_6_0_t1130;
    FSM_fft_64_stage_6_0_t1139[FSM_fft_64_stage_6_0_t1132 * 32 +: 32] = FSM_fft_64_stage_6_0_t1135 - FSM_fft_64_stage_6_0_t1138;
    FSM_fft_64_stage_6_0_t1140 = 32'b00000000000000000000000000011001;
    FSM_fft_64_stage_6_0_t1141 = FSM_fft_64_stage_6_0_t1140[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1142 = 32'b00000000000000000000000000011001;
    FSM_fft_64_stage_6_0_t1143 = FSM_fft_64_stage_6_0_t1142[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1144 = i_data_in_imag[FSM_fft_64_stage_6_0_t1143 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1145 = 32'b00000000000000000000000000111001;
    FSM_fft_64_stage_6_0_t1146 = FSM_fft_64_stage_6_0_t1145[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1147 = i_data_in_imag[FSM_fft_64_stage_6_0_t1146 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1148 = FSM_fft_64_stage_6_0_t1144 + FSM_fft_64_stage_6_0_t1147;
    FSM_fft_64_stage_6_0_t1149 = FSM_fft_64_stage_6_0_t1148[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t1150 = FSM_fft_64_stage_6_0_t1139;
    FSM_fft_64_stage_6_0_t1150[FSM_fft_64_stage_6_0_t1141 * 32 +: 32] = FSM_fft_64_stage_6_0_t1149;
    FSM_fft_64_stage_6_0_t1151 = 32'b00000000000000000000000000111001;
    FSM_fft_64_stage_6_0_t1152 = FSM_fft_64_stage_6_0_t1151[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1153 = 32'b00000000000000000000000000011001;
    FSM_fft_64_stage_6_0_t1154 = FSM_fft_64_stage_6_0_t1153[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1155 = i_data_in_imag[FSM_fft_64_stage_6_0_t1154 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1156 = 32'b00000000000000000000000000111001;
    FSM_fft_64_stage_6_0_t1157 = FSM_fft_64_stage_6_0_t1156[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1158 = i_data_in_imag[FSM_fft_64_stage_6_0_t1157 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1159 = FSM_fft_64_stage_6_0_t1150;
    FSM_fft_64_stage_6_0_t1159[FSM_fft_64_stage_6_0_t1152 * 32 +: 32] = FSM_fft_64_stage_6_0_t1155 - FSM_fft_64_stage_6_0_t1158;
    FSM_fft_64_stage_6_0_t1160 = 32'b00000000000000000000000000011010;
    FSM_fft_64_stage_6_0_t1161 = FSM_fft_64_stage_6_0_t1160[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1162 = 32'b00000000000000000000000000011010;
    FSM_fft_64_stage_6_0_t1163 = FSM_fft_64_stage_6_0_t1162[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1164 = i_data_in_imag[FSM_fft_64_stage_6_0_t1163 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1165 = 32'b00000000000000000000000000111010;
    FSM_fft_64_stage_6_0_t1166 = FSM_fft_64_stage_6_0_t1165[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1167 = i_data_in_imag[FSM_fft_64_stage_6_0_t1166 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1168 = FSM_fft_64_stage_6_0_t1164 + FSM_fft_64_stage_6_0_t1167;
    FSM_fft_64_stage_6_0_t1169 = FSM_fft_64_stage_6_0_t1168[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t1170 = FSM_fft_64_stage_6_0_t1159;
    FSM_fft_64_stage_6_0_t1170[FSM_fft_64_stage_6_0_t1161 * 32 +: 32] = FSM_fft_64_stage_6_0_t1169;
    FSM_fft_64_stage_6_0_t1171 = 32'b00000000000000000000000000111010;
    FSM_fft_64_stage_6_0_t1172 = FSM_fft_64_stage_6_0_t1171[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1173 = 32'b00000000000000000000000000011010;
    FSM_fft_64_stage_6_0_t1174 = FSM_fft_64_stage_6_0_t1173[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1175 = i_data_in_imag[FSM_fft_64_stage_6_0_t1174 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1176 = 32'b00000000000000000000000000111010;
    FSM_fft_64_stage_6_0_t1177 = FSM_fft_64_stage_6_0_t1176[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1178 = i_data_in_imag[FSM_fft_64_stage_6_0_t1177 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1179 = FSM_fft_64_stage_6_0_t1170;
    FSM_fft_64_stage_6_0_t1179[FSM_fft_64_stage_6_0_t1172 * 32 +: 32] = FSM_fft_64_stage_6_0_t1175 - FSM_fft_64_stage_6_0_t1178;
    FSM_fft_64_stage_6_0_t1180 = 32'b00000000000000000000000000011011;
    FSM_fft_64_stage_6_0_t1181 = FSM_fft_64_stage_6_0_t1180[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1182 = 32'b00000000000000000000000000011011;
    FSM_fft_64_stage_6_0_t1183 = FSM_fft_64_stage_6_0_t1182[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1184 = i_data_in_imag[FSM_fft_64_stage_6_0_t1183 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1185 = 32'b00000000000000000000000000111011;
    FSM_fft_64_stage_6_0_t1186 = FSM_fft_64_stage_6_0_t1185[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1187 = i_data_in_imag[FSM_fft_64_stage_6_0_t1186 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1188 = FSM_fft_64_stage_6_0_t1184 + FSM_fft_64_stage_6_0_t1187;
    FSM_fft_64_stage_6_0_t1189 = FSM_fft_64_stage_6_0_t1188[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t1190 = FSM_fft_64_stage_6_0_t1179;
    FSM_fft_64_stage_6_0_t1190[FSM_fft_64_stage_6_0_t1181 * 32 +: 32] = FSM_fft_64_stage_6_0_t1189;
    FSM_fft_64_stage_6_0_t1191 = 32'b00000000000000000000000000111011;
    FSM_fft_64_stage_6_0_t1192 = FSM_fft_64_stage_6_0_t1191[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1193 = 32'b00000000000000000000000000011011;
    FSM_fft_64_stage_6_0_t1194 = FSM_fft_64_stage_6_0_t1193[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1195 = i_data_in_imag[FSM_fft_64_stage_6_0_t1194 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1196 = 32'b00000000000000000000000000111011;
    FSM_fft_64_stage_6_0_t1197 = FSM_fft_64_stage_6_0_t1196[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1198 = i_data_in_imag[FSM_fft_64_stage_6_0_t1197 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1199 = FSM_fft_64_stage_6_0_t1190;
    FSM_fft_64_stage_6_0_t1199[FSM_fft_64_stage_6_0_t1192 * 32 +: 32] = FSM_fft_64_stage_6_0_t1195 - FSM_fft_64_stage_6_0_t1198;
    FSM_fft_64_stage_6_0_t1200 = 32'b00000000000000000000000000011100;
    FSM_fft_64_stage_6_0_t1201 = FSM_fft_64_stage_6_0_t1200[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1202 = 32'b00000000000000000000000000011100;
    FSM_fft_64_stage_6_0_t1203 = FSM_fft_64_stage_6_0_t1202[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1204 = i_data_in_imag[FSM_fft_64_stage_6_0_t1203 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1205 = 32'b00000000000000000000000000111100;
    FSM_fft_64_stage_6_0_t1206 = FSM_fft_64_stage_6_0_t1205[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1207 = i_data_in_imag[FSM_fft_64_stage_6_0_t1206 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1208 = FSM_fft_64_stage_6_0_t1204 + FSM_fft_64_stage_6_0_t1207;
    FSM_fft_64_stage_6_0_t1209 = FSM_fft_64_stage_6_0_t1208[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t1210 = FSM_fft_64_stage_6_0_t1199;
    FSM_fft_64_stage_6_0_t1210[FSM_fft_64_stage_6_0_t1201 * 32 +: 32] = FSM_fft_64_stage_6_0_t1209;
    FSM_fft_64_stage_6_0_t1211 = 32'b00000000000000000000000000111100;
    FSM_fft_64_stage_6_0_t1212 = FSM_fft_64_stage_6_0_t1211[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1213 = 32'b00000000000000000000000000011100;
    FSM_fft_64_stage_6_0_t1214 = FSM_fft_64_stage_6_0_t1213[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1215 = i_data_in_imag[FSM_fft_64_stage_6_0_t1214 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1216 = 32'b00000000000000000000000000111100;
    FSM_fft_64_stage_6_0_t1217 = FSM_fft_64_stage_6_0_t1216[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1218 = i_data_in_imag[FSM_fft_64_stage_6_0_t1217 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1219 = FSM_fft_64_stage_6_0_t1210;
    FSM_fft_64_stage_6_0_t1219[FSM_fft_64_stage_6_0_t1212 * 32 +: 32] = FSM_fft_64_stage_6_0_t1215 - FSM_fft_64_stage_6_0_t1218;
    FSM_fft_64_stage_6_0_t1220 = 32'b00000000000000000000000000011101;
    FSM_fft_64_stage_6_0_t1221 = FSM_fft_64_stage_6_0_t1220[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1222 = 32'b00000000000000000000000000011101;
    FSM_fft_64_stage_6_0_t1223 = FSM_fft_64_stage_6_0_t1222[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1224 = i_data_in_imag[FSM_fft_64_stage_6_0_t1223 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1225 = 32'b00000000000000000000000000111101;
    FSM_fft_64_stage_6_0_t1226 = FSM_fft_64_stage_6_0_t1225[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1227 = i_data_in_imag[FSM_fft_64_stage_6_0_t1226 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1228 = FSM_fft_64_stage_6_0_t1224 + FSM_fft_64_stage_6_0_t1227;
    FSM_fft_64_stage_6_0_t1229 = FSM_fft_64_stage_6_0_t1228[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t1230 = FSM_fft_64_stage_6_0_t1219;
    FSM_fft_64_stage_6_0_t1230[FSM_fft_64_stage_6_0_t1221 * 32 +: 32] = FSM_fft_64_stage_6_0_t1229;
    FSM_fft_64_stage_6_0_t1231 = 32'b00000000000000000000000000111101;
    FSM_fft_64_stage_6_0_t1232 = FSM_fft_64_stage_6_0_t1231[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1233 = 32'b00000000000000000000000000011101;
    FSM_fft_64_stage_6_0_t1234 = FSM_fft_64_stage_6_0_t1233[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1235 = i_data_in_imag[FSM_fft_64_stage_6_0_t1234 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1236 = 32'b00000000000000000000000000111101;
    FSM_fft_64_stage_6_0_t1237 = FSM_fft_64_stage_6_0_t1236[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1238 = i_data_in_imag[FSM_fft_64_stage_6_0_t1237 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1239 = FSM_fft_64_stage_6_0_t1230;
    FSM_fft_64_stage_6_0_t1239[FSM_fft_64_stage_6_0_t1232 * 32 +: 32] = FSM_fft_64_stage_6_0_t1235 - FSM_fft_64_stage_6_0_t1238;
    FSM_fft_64_stage_6_0_t1240 = 32'b00000000000000000000000000011110;
    FSM_fft_64_stage_6_0_t1241 = FSM_fft_64_stage_6_0_t1240[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1242 = 32'b00000000000000000000000000011110;
    FSM_fft_64_stage_6_0_t1243 = FSM_fft_64_stage_6_0_t1242[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1244 = i_data_in_imag[FSM_fft_64_stage_6_0_t1243 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1245 = 32'b00000000000000000000000000111110;
    FSM_fft_64_stage_6_0_t1246 = FSM_fft_64_stage_6_0_t1245[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1247 = i_data_in_imag[FSM_fft_64_stage_6_0_t1246 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1248 = FSM_fft_64_stage_6_0_t1244 + FSM_fft_64_stage_6_0_t1247;
    FSM_fft_64_stage_6_0_t1249 = FSM_fft_64_stage_6_0_t1248[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t1250 = FSM_fft_64_stage_6_0_t1239;
    FSM_fft_64_stage_6_0_t1250[FSM_fft_64_stage_6_0_t1241 * 32 +: 32] = FSM_fft_64_stage_6_0_t1249;
    FSM_fft_64_stage_6_0_t1251 = 32'b00000000000000000000000000111110;
    FSM_fft_64_stage_6_0_t1252 = FSM_fft_64_stage_6_0_t1251[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1253 = 32'b00000000000000000000000000011110;
    FSM_fft_64_stage_6_0_t1254 = FSM_fft_64_stage_6_0_t1253[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1255 = i_data_in_imag[FSM_fft_64_stage_6_0_t1254 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1256 = 32'b00000000000000000000000000111110;
    FSM_fft_64_stage_6_0_t1257 = FSM_fft_64_stage_6_0_t1256[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1258 = i_data_in_imag[FSM_fft_64_stage_6_0_t1257 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1259 = FSM_fft_64_stage_6_0_t1250;
    FSM_fft_64_stage_6_0_t1259[FSM_fft_64_stage_6_0_t1252 * 32 +: 32] = FSM_fft_64_stage_6_0_t1255 - FSM_fft_64_stage_6_0_t1258;
    FSM_fft_64_stage_6_0_t1260 = 32'b00000000000000000000000000011111;
    FSM_fft_64_stage_6_0_t1261 = FSM_fft_64_stage_6_0_t1260[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1262 = 32'b00000000000000000000000000011111;
    FSM_fft_64_stage_6_0_t1263 = FSM_fft_64_stage_6_0_t1262[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1264 = i_data_in_imag[FSM_fft_64_stage_6_0_t1263 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1265 = 32'b00000000000000000000000000111111;
    FSM_fft_64_stage_6_0_t1266 = FSM_fft_64_stage_6_0_t1265[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1267 = i_data_in_imag[FSM_fft_64_stage_6_0_t1266 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1268 = FSM_fft_64_stage_6_0_t1264 + FSM_fft_64_stage_6_0_t1267;
    FSM_fft_64_stage_6_0_t1269 = FSM_fft_64_stage_6_0_t1268[6'b0 * 1 +: 32 * 1];
    FSM_fft_64_stage_6_0_t1270 = FSM_fft_64_stage_6_0_t1259;
    FSM_fft_64_stage_6_0_t1270[FSM_fft_64_stage_6_0_t1261 * 32 +: 32] = FSM_fft_64_stage_6_0_t1269;
    FSM_fft_64_stage_6_0_t1271 = 32'b00000000000000000000000000111111;
    FSM_fft_64_stage_6_0_t1272 = FSM_fft_64_stage_6_0_t1271[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1273 = 32'b00000000000000000000000000011111;
    FSM_fft_64_stage_6_0_t1274 = FSM_fft_64_stage_6_0_t1273[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1275 = i_data_in_imag[FSM_fft_64_stage_6_0_t1274 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1276 = 32'b00000000000000000000000000111111;
    FSM_fft_64_stage_6_0_t1277 = FSM_fft_64_stage_6_0_t1276[5'b0 * 1 +: 6 * 1];
    FSM_fft_64_stage_6_0_t1278 = i_data_in_imag[FSM_fft_64_stage_6_0_t1277 * 32 +: 32];
    FSM_fft_64_stage_6_0_t1279 = FSM_fft_64_stage_6_0_t1270;
    FSM_fft_64_stage_6_0_t1279[FSM_fft_64_stage_6_0_t1272 * 32 +: 32] = FSM_fft_64_stage_6_0_t1275 - FSM_fft_64_stage_6_0_t1278;
end

assign FSM_fft_64_stage_6_0_in_ready = 1'b1;

always @(posedge clk) begin
    FSM_fft_64_stage_6_0_st_dummy_reg <= FSM_fft_64_stage_6_0_st_dummy_reg;
    if (rst) begin
        FSM_fft_64_stage_6_0_st_dummy_reg <= 32'b0;
    end
end
/* End submodules of fft_64_stage_6 */
/* End module fft_64_stage_6 */
endgenerate
endmodule
